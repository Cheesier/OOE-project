library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity alu is
    Port (  clk : in STD_LOGIC;
            op : in STD_LOGIC_VECTOR(3 downto 0);
            A, B : in STD_LOGIC_VECTOR(15 downto 0);
            result : out STD_LOGIC_VECTOR(15 downto 0);
            carry, zero, negative, overflow : out STD_LOGIC);
end alu;

architecture alu_one of alu is
    signal value : STD_LOGIC_VECTOR(16 downto 0) := "00000000000000000";
    signal useflag : STD_LOGIC := '0';

begin
    process(A, B, op) begin
        case op is
            when "0001" => value <= '0' & B; --databus
                           useflag <= '1';
            when "0011" => value <= "00000000000000000"; --nollställ
                           useflag <= '1';
            when "0100" => value <= STD_LOGIC_VECTOR('0' & unsigned(A) + unsigned(B)); --add
                           useflag <= '1';
            when "0101" => value <= ('0' & A) - B; --sub
                           useflag <= '1';
            when "0110" => value <= '0' & A and '0' & B; -- and
                           useflag <= '1';
            when "0111" => value <= '0' & A or '0' & B; -- or
                           useflag <= '1';
            when "1000" => value <= STD_LOGIC_VECTOR('0' & unsigned(A) + unsigned(B)); --add noflag
                           useflag <= '0';
            when "1001" => value <= a & '0'; -- ASL/LSL
                           useflag <= '1';
            when "1011" => value <= a(0) & a(15) & a(15 downto 1); -- ASR
                           useflag <= '1';
            when "1101" => value <= a(0) & '0' & a(15 downto 1); -- LSR
                           useflag <= '1';
            when others => value <= '0' & A; -- AR
                           useflag <= '0';
        end case;
    end process;
    
    process(clk) begin
    --process(value, useflag) begin
        if rising_edge(clk) then
            result <= value(15 downto 0);
            if useflag = '1' then
                if value(15 downto 0) = X"0000" then
                    zero <= '1';
                else
                    zero <= '0';
                end if;
                if value(16) = '1' then carry <= '1';
                else carry <= '0'; 
                end if;
                if value(15) = '1' then negative <= '1'; 
                else negative <= '0'; 
                end if;
                if value(16) /= value(15) then overflow <= '1';
                else overflow <= '0';
                end if;
            end if; 
        end if;
    end process;
end alu_one;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity cpu is
    Port (clk,rst : in  STD_LOGIC;
        sw: in STD_LOGIC_VECTOR(7 downto 0);
        seg: out  STD_LOGIC_VECTOR(7 downto 0);
        an : out  STD_LOGIC_VECTOR (3 downto 0);
        led : out STD_LOGIC_VECTOR (7 downto 0);
        vr_we : out STD_LOGIC;
        vr_addr : out STD_LOGIC_VECTOR(4 downto 0);
        vr_i : out STD_LOGIC_VECTOR(15 downto 0);
        vr_o : in STD_LOGIC_VECTOR(15 downto 0);
        fV: in STD_LOGIC;
        up, right, down, left : in STD_LOGIC);
end cpu;

architecture cpu_one of cpu is

    component leddriver
        Port ( clk,rst : in  STD_LOGIC;
           seg : out  STD_LOGIC_VECTOR(7 downto 0);
           an : out  STD_LOGIC_VECTOR (3 downto 0);
           led : out STD_LOGIC_VECTOR (7 downto 0);
           value : in  STD_LOGIC_VECTOR (15 downto 0);
           ledval : in STD_LOGIC_VECTOR (7 downto 0));
    end component;

    component alu
        Port (clk : in STD_LOGIC;
            op : in STD_LOGIC_VECTOR(3 downto 0);
            A, B : in STD_LOGIC_VECTOR(15 downto 0);
            result : out STD_LOGIC_VECTOR(15 downto 0);
            carry, zero, negative, overflow : out STD_LOGIC);
    end component;

    signal databus : STD_LOGIC_VECTOR(15 downto 0) := X"0000";

    -- Registers
    signal rASR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rIR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rPC : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rDR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rAR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rHR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rSP : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rLC : STD_LOGIC_VECTOR(7 downto 0) := X"00";

    -- Flags
    signal fZ : STD_LOGIC := '1';
    signal fN : STD_LOGIC := '0';
    signal fC : STD_LOGIC := '0';
    signal fO : STD_LOGIC := '0';
    signal fL : STD_LOGIC := '0';

    -- Primary memory
    type PrimMem_type is array (0 to 2047) of STD_LOGIC_VECTOR(15 downto 0);
    signal PrimMem : PrimMem_type := (  0=> X"0100",1=> X"0000",2=> X"0110",3=> X"00d0",4=> X"0140",5=> X"00f0",6=> X"0120",7=> X"0001",8=> X"0130",9=> X"0002",10=> X"0540",11=> X"0022",12=> X"0510",13=> X"0023",14=> X"0500",15=> X"0024",16=> X"0500",17=> X"0025",18=> X"0500",19=> X"0026",20=> X"0500",21=> X"0027",22=> X"0500",23=> X"0028",24=> X"0500",25=> X"002d",26=> X"0500",27=> X"002e",28=> X"0520",29=> X"002f",30=> X"0530",31=> X"0030",32=> X"0d00",33=> X"003f",34=> X"0000",35=> X"0000",36=> X"0000",37=> X"0000",38=> X"0000",39=> X"0000",40=> X"0000",41=> X"0000",42=> X"0000",43=> X"0000",44=> X"0000",45=> X"0000",46=> X"0000",47=> X"0000",48=> X"0000",49=> X"0000",50=> X"0000",51=> X"0000",52=> X"0000",53=> X"0000",54=> X"0002",55=> X"0000",56=> X"0000",57=> X"0000",58=> X"fffc",59=> X"0000",60=> X"0000",61=> X"0640",62=> X"03c0",63=> X"3500",64=> X"07ff",65=> X"2500",66=> X"0064",67=> X"2500",68=> X"00b9",69=> X"2500",70=> X"00f0",71=> X"2500",72=> X"012d",73=> X"2500",74=> X"014c",75=> X"0200",76=> X"0022",77=> X"4500",78=> X"0fff",79=> X"0500",80=> X"0022",81=> X"2500",82=> X"016b",83=> X"2500",84=> X"01d8",85=> X"2500",86=> X"0309",87=> X"2500",88=> X"031c",89=> X"0220",90=> X"0022",91=> X"0230",92=> X"0022",93=> X"0240",94=> X"002d",95=> X"0250",96=> X"0025",97=> X"1c00",98=> X"0d00",99=> X"0041",100=> X"2d00",101=> X"0000",102=> X"2d10",103=> X"0000",104=> X"0200",105=> X"8004",106=> X"4500",107=> X"0001",108=> X"0500",109=> X"0024",110=> X"0200",111=> X"8000",112=> X"0210",113=> X"0033",114=> X"4a10",115=> X"0034",116=> X"0801",117=> X"2100",118=> X"0002",119=> X"1900",120=> X"0081",121=> X"0100",122=> X"0020",123=> X"0500",124=> X"0028",125=> X"0100",126=> X"0000",127=> X"0500",128=> X"0027",129=> X"0200",130=> X"8001",131=> X"0210",132=> X"8003",133=> X"2001",134=> X"4d00",135=> X"0094",136=> X"1500",137=> X"009e",138=> X"0110",139=> X"0002",140=> X"0510",141=> X"002e",142=> X"0110",143=> X"0001",144=> X"0510",145=> X"002d",146=> X"0d00",147=> X"00b4",148=> X"0110",149=> X"0002",150=> X"0510",151=> X"002e",152=> X"0110",153=> X"0000",154=> X"0510",155=> X"002d",156=> X"0d00",157=> X"00b4",158=> X"0210",159=> X"0026",160=> X"2110",161=> X"0000",162=> X"1500",163=> X"00b0",164=> X"5610",165=> X"0025",166=> X"0910",167=> X"0001",168=> X"0510",169=> X"002d",170=> X"0110",171=> X"0001",172=> X"0510",173=> X"002e",174=> X"0d00",175=> X"00b4",176=> X"0110",177=> X"0000",178=> X"0510",179=> X"002e",180=> X"3110",181=> X"0000",182=> X"3100",183=> X"0000",184=> X"2800",185=> X"2d00",186=> X"0000",187=> X"2d10",188=> X"0000",189=> X"0200",190=> X"0025",191=> X"2200",192=> X"002d",193=> X"1500",194=> X"00c5",195=> X"1900",196=> X"00cd",197=> X"0200",198=> X"0026",199=> X"0a00",200=> X"002e",201=> X"0500",202=> X"0026",203=> X"0d00",204=> X"00e1",205=> X"0200",206=> X"0026",207=> X"3a00",208=> X"002e",209=> X"4d00",210=> X"00d7",211=> X"0500",212=> X"0026",213=> X"0d00",214=> X"00e1",215=> X"5600",216=> X"0026",217=> X"0500",218=> X"0026",219=> X"5600",220=> X"0025",221=> X"0900",222=> X"0001",223=> X"0500",224=> X"0025",225=> X"0200",226=> X"0026",227=> X"2100",228=> X"0018",229=> X"4d00",230=> X"00eb",231=> X"0100",232=> X"0018",233=> X"0500",234=> X"0026",235=> X"3110",236=> X"0000",237=> X"3100",238=> X"0000",239=> X"2800",240=> X"2d00",241=> X"0000",242=> X"2d10",243=> X"0000",244=> X"0200",245=> X"0027",246=> X"2200",247=> X"002f",248=> X"1500",249=> X"00fc",250=> X"1900",251=> X"0104",252=> X"0200",253=> X"0028",254=> X"0a00",255=> X"0030",256=> X"0500",257=> X"0028",258=> X"0d00",259=> X"0118",260=> X"0200",261=> X"0028",262=> X"3a00",263=> X"0030",264=> X"4d00",265=> X"010e",266=> X"0500",267=> X"0028",268=> X"0d00",269=> X"0118",270=> X"5600",271=> X"0028",272=> X"0500",273=> X"0028",274=> X"5600",275=> X"0027",276=> X"0900",277=> X"0001",278=> X"0500",279=> X"0027",280=> X"0200",281=> X"0027",282=> X"2100",283=> X"0001",284=> X"1900",285=> X"0128",286=> X"0200",287=> X"0028",288=> X"2100",289=> X"0020",290=> X"4d00",291=> X"0128",292=> X"0100",293=> X"0020",294=> X"0500",295=> X"0028",296=> X"3110",297=> X"0000",298=> X"3100",299=> X"0000",300=> X"2800",301=> X"2d00",302=> X"0000",303=> X"2d10",304=> X"0000",305=> X"2d80",306=> X"0000",307=> X"0200",308=> X"0026",309=> X"0210",310=> X"0022",311=> X"3d00",312=> X"0003",313=> X"0280",314=> X"0025",315=> X"2180",316=> X"0001",317=> X"1900",318=> X"0142",319=> X"0810",320=> X"0d00",321=> X"0143",322=> X"3810",323=> X"0510",324=> X"0022",325=> X"3180",326=> X"0000",327=> X"3110",328=> X"0000",329=> X"3100",330=> X"0000",331=> X"2800",332=> X"2d00",333=> X"0000",334=> X"2d10",335=> X"0000",336=> X"2d80",337=> X"0000",338=> X"0200",339=> X"0028",340=> X"0210",341=> X"0023",342=> X"3d00",343=> X"0003",344=> X"0280",345=> X"0027",346=> X"2180",347=> X"0001",348=> X"1900",349=> X"0161",350=> X"0810",351=> X"0d00",352=> X"0162",353=> X"3810",354=> X"0510",355=> X"0023",356=> X"3180",357=> X"0000",358=> X"3110",359=> X"0000",360=> X"3100",361=> X"0000",362=> X"2800",363=> X"2d00",364=> X"0000",365=> X"2d10",366=> X"0000",367=> X"2d20",368=> X"0000",369=> X"0200",370=> X"0022",371=> X"0210",372=> X"0023",373=> X"2500",374=> X"01a0",375=> X"0500",376=> X"0031",377=> X"0200",378=> X"0022",379=> X"0900",380=> X"000f",381=> X"0210",382=> X"0023",383=> X"2500",384=> X"01a0",385=> X"0500",386=> X"0032",387=> X"0200",388=> X"0022",389=> X"0210",390=> X"0023",391=> X"0910",392=> X"000f",393=> X"2500",394=> X"01a0",395=> X"0500",396=> X"0033",397=> X"0200",398=> X"0022",399=> X"0900",400=> X"000f",401=> X"0210",402=> X"0023",403=> X"0910",404=> X"000f",405=> X"2500",406=> X"01a0",407=> X"0500",408=> X"0034",409=> X"3120",410=> X"0000",411=> X"3110",412=> X"0000",413=> X"3100",414=> X"0000",415=> X"2800",416=> X"2d20",417=> X"0000",418=> X"2d30",419=> X"0000",420=> X"2d40",421=> X"0000",422=> X"2df0",423=> X"0000",424=> X"3d00",425=> X"0004",426=> X"3d10",427=> X"0004",428=> X"0050",429=> X"3d00",430=> X"0004",431=> X"4500",432=> X"0007",433=> X"4110",434=> X"0003",435=> X"0801",436=> X"02f0",437=> X"0024",438=> X"03ff",439=> X"003d",440=> X"08f0",441=> X"032f",442=> X"0000",443=> X"0005",444=> X"4500",445=> X"000f",446=> X"0130",447=> X"000f",448=> X"3830",449=> X"0140",450=> X"0001",451=> X"4043",452=> X"4424",453=> X"2120",454=> X"0000",455=> X"1500",456=> X"01cd",457=> X"0100",458=> X"0001",459=> X"0d00",460=> X"01cf",461=> X"0100",462=> X"0000",463=> X"31f0",464=> X"0000",465=> X"3140",466=> X"0000",467=> X"3130",468=> X"0000",469=> X"3120",470=> X"0000",471=> X"2800",472=> X"2d00",473=> X"0000",474=> X"2d10",475=> X"0000",476=> X"2d20",477=> X"0000",478=> X"0200",479=> X"0031",480=> X"2100",481=> X"0001",482=> X"1500",483=> X"01f8",484=> X"0200",485=> X"0032",486=> X"2100",487=> X"0001",488=> X"1500",489=> X"0206",490=> X"0200",491=> X"0033",492=> X"2100",493=> X"0001",494=> X"1500",495=> X"020e",496=> X"0200",497=> X"0034",498=> X"2100",499=> X"0001",500=> X"1500",501=> X"02fe",502=> X"0d00",503=> X"0302",504=> X"0200",505=> X"0032",506=> X"2100",507=> X"0001",508=> X"1500",509=> X"0216",510=> X"0200",511=> X"0033",512=> X"2100",513=> X"0001",514=> X"1500",515=> X"0234",516=> X"0d00",517=> X"02dc",518=> X"0200",519=> X"0034",520=> X"2100",521=> X"0001",522=> X"1500",523=> X"024c",524=> X"0d00",525=> X"02ee",526=> X"0200",527=> X"0034",528=> X"2100",529=> X"0001",530=> X"1500",531=> X"0261",532=> X"0d00",533=> X"02fc",534=> X"0100",535=> X"0000",536=> X"0600",537=> X"0028",538=> X"0200",539=> X"0033",540=> X"2100",541=> X"0001",542=> X"1500",543=> X"0270",544=> X"0200",545=> X"0034",546=> X"2100",547=> X"0001",548=> X"1500",549=> X"028e",550=> X"0210",551=> X"0023",552=> X"4510",553=> X"000f",554=> X"0220",555=> X"0023",556=> X"0130",557=> X"0010",558=> X"3831",559=> X"0823",560=> X"0520",561=> X"0023",562=> X"0d00",563=> X"0302",564=> X"0100",565=> X"0000",566=> X"0600",567=> X"0026",568=> X"0200",569=> X"0034",570=> X"2100",571=> X"0001",572=> X"1500",573=> X"02a9",574=> X"0210",575=> X"0022",576=> X"4510",577=> X"000f",578=> X"0220",579=> X"0022",580=> X"0130",581=> X"0010",582=> X"3831",583=> X"0823",584=> X"0520",585=> X"0022",586=> X"0d00",587=> X"0302",588=> X"0100",589=> X"0000",590=> X"0600",591=> X"0026",592=> X"0200",593=> X"0033",594=> X"2100",595=> X"0001",596=> X"1500",597=> X"02c4",598=> X"0210",599=> X"0022",600=> X"4510",601=> X"000f",602=> X"0220",603=> X"0022",604=> X"3821",605=> X"0520",606=> X"0022",607=> X"0d00",608=> X"0302",609=> X"0100",610=> X"0000",611=> X"0600",612=> X"0028",613=> X"0210",614=> X"0023",615=> X"4510",616=> X"000f",617=> X"0220",618=> X"0023",619=> X"3821",620=> X"0520",621=> X"0023",622=> X"0d00",623=> X"0302",624=> X"0210",625=> X"0023",626=> X"4510",627=> X"000f",628=> X"0220",629=> X"0023",630=> X"0130",631=> X"0010",632=> X"3831",633=> X"0823",634=> X"0520",635=> X"0023",636=> X"0100",637=> X"0000",638=> X"0600",639=> X"0026",640=> X"0210",641=> X"0022",642=> X"4510",643=> X"000f",644=> X"0220",645=> X"0022",646=> X"0130",647=> X"0010",648=> X"3831",649=> X"0823",650=> X"0520",651=> X"0022",652=> X"0d00",653=> X"0302",654=> X"0210",655=> X"0023",656=> X"4510",657=> X"000f",658=> X"0220",659=> X"0023",660=> X"0130",661=> X"0010",662=> X"3831",663=> X"0823",664=> X"0520",665=> X"0023",666=> X"0100",667=> X"0000",668=> X"0600",669=> X"0026",670=> X"0210",671=> X"0022",672=> X"4510",673=> X"000f",674=> X"0220",675=> X"0022",676=> X"3821",677=> X"0520",678=> X"0022",679=> X"0d00",680=> X"0302",681=> X"0210",682=> X"0022",683=> X"4510",684=> X"000f",685=> X"0220",686=> X"0022",687=> X"0130",688=> X"0010",689=> X"3831",690=> X"0823",691=> X"0520",692=> X"0022",693=> X"0100",694=> X"0000",695=> X"0600",696=> X"0028",697=> X"0210",698=> X"0023",699=> X"4510",700=> X"000f",701=> X"0220",702=> X"0023",703=> X"3821",704=> X"0520",705=> X"0023",706=> X"0d00",707=> X"0302",708=> X"0210",709=> X"0022",710=> X"4510",711=> X"000f",712=> X"0220",713=> X"0022",714=> X"3821",715=> X"0520",716=> X"0022",717=> X"0100",718=> X"0000",719=> X"0600",720=> X"0028",721=> X"0210",722=> X"0023",723=> X"4510",724=> X"000f",725=> X"0220",726=> X"0023",727=> X"3821",728=> X"0520",729=> X"0023",730=> X"0d00",731=> X"0302",732=> X"0100",733=> X"0000",734=> X"0600",735=> X"0028",736=> X"0210",737=> X"0023",738=> X"4510",739=> X"000f",740=> X"0220",741=> X"0023",742=> X"0130",743=> X"0010",744=> X"3831",745=> X"0823",746=> X"0520",747=> X"0023",748=> X"0d00",749=> X"0302",750=> X"0210",751=> X"0023",752=> X"4510",753=> X"000f",754=> X"0220",755=> X"0023",756=> X"0130",757=> X"0010",758=> X"3831",759=> X"0823",760=> X"0520",761=> X"0023",762=> X"0d00",763=> X"0302",764=> X"0d00",765=> X"0261",766=> X"0d00",767=> X"0261",768=> X"0d00",769=> X"0302",770=> X"3120",771=> X"0000",772=> X"3110",773=> X"0000",774=> X"3100",775=> X"0000",776=> X"2800",777=> X"2d00",778=> X"0000",779=> X"0200",780=> X"0022",781=> X"3d00",782=> X"0003",783=> X"5400",784=> X"0500",785=> X"0037",786=> X"0200",787=> X"0022",788=> X"3d00",789=> X"0004",790=> X"5400",791=> X"0500",792=> X"0038",793=> X"3100",794=> X"0000",795=> X"2800",796=> X"2d00",797=> X"0000",798=> X"02f0",799=> X"0024",800=> X"0200",801=> X"0022",802=> X"0b0f",803=> X"0035",804=> X"0500",805=> X"9000",806=> X"0200",807=> X"0023",808=> X"0b0f",809=> X"0039",810=> X"0500",811=> X"9001",812=> X"0200",813=> X"0035",814=> X"0500",815=> X"9010",816=> X"0200",817=> X"0039",818=> X"0500",819=> X"9011",820=> X"0200",821=> X"0036",822=> X"0500",823=> X"9012",824=> X"0200",825=> X"003a",826=> X"0500",827=> X"9013",828=> X"0200",829=> X"0037",830=> X"0500",831=> X"9014",832=> X"0200",833=> X"003b",834=> X"0500",835=> X"9015",836=> X"0200",837=> X"0038",838=> X"0500",839=> X"9016",840=> X"0200",841=> X"003c",842=> X"0500",843=> X"9017",844=> X"0200",845=> X"0024",846=> X"4100",847=> X"000e",848=> X"0500",849=> X"901a",850=> X"3100",851=> X"0000",852=> X"2800",853=> X"2d00",854=> X"0000",855=> X"0200",856=> X"0023",857=> X"3a00",858=> X"8000",859=> X"0a00",860=> X"8002",861=> X"0500",862=> X"0023",863=> X"0200",864=> X"0022",865=> X"0a00",866=> X"8001",867=> X"3a00",868=> X"8003",869=> X"0500",870=> X"0022",871=> X"3100",872=> X"0000",873=> X"2800",
                                        960=> X"ffff",961=> X"ffff",962=> X"ff00",963=> X"0000",964=> X"0000",965=> X"0000",966=> X"0000",967=> X"0000",968=> X"8000",969=> X"0000",970=> X"0100",971=> X"0000",972=> X"0000",973=> X"0000",974=> X"0000",975=> X"0000",976=> X"8000",977=> X"0000",978=> X"0100",979=> X"0000",980=> X"0000",981=> X"0000",982=> X"0000",983=> X"0000",984=> X"8000",985=> X"0000",986=> X"0100",987=> X"0000",988=> X"0000",989=> X"0000",990=> X"0000",991=> X"0000",992=> X"8007",993=> X"0000",994=> X"0100",995=> X"0000",996=> X"0000",997=> X"0000",998=> X"0000",999=> X"0000",1000=> X"8008",1001=> X"8000",1002=> X"0100",1003=> X"0000",1004=> X"0000",1005=> X"0000",1006=> X"0000",1007=> X"0000",1008=> X"8010",1009=> X"4000",1010=> X"0100",1011=> X"0000",1012=> X"0000",1013=> X"0000",1014=> X"0000",1015=> X"0000",1016=> X"8010",1017=> X"4000",1018=> X"0100",1019=> X"0000",1020=> X"0000",1021=> X"0000",1022=> X"0000",1023=> X"0000",1024=> X"8020",1025=> X"2000",1026=> X"0100",1027=> X"0000",1028=> X"0000",1029=> X"0000",1030=> X"0000",1031=> X"0000",1032=> X"8020",1033=> X"3c00",1034=> X"0100",1035=> X"0000",1036=> X"0000",1037=> X"0000",1038=> X"0000",1039=> X"0000",1040=> X"8020",1041=> X"2000",1042=> X"0100",1043=> X"0000",1044=> X"0000",1045=> X"0000",1046=> X"0000",1047=> X"0000",1048=> X"8020",1049=> X"2000",1050=> X"1d00",1051=> X"0000",1052=> X"0000",1053=> X"0000",1054=> X"0000",1055=> X"0000",1056=> X"8020",1057=> X"2000",1058=> X"1100",1059=> X"0000",1060=> X"0000",1061=> X"0000",1062=> X"0000",1063=> X"0000",1064=> X"8000",1065=> X"03ff",1066=> X"f100",1067=> X"0000",1068=> X"0000",1069=> X"0000",1070=> X"0000",1071=> X"0000",1072=> X"8000",1073=> X"0200",1074=> X"1100",1075=> X"0000",1076=> X"0000",1077=> X"0000",1078=> X"0000",1079=> X"0000",1080=> X"e000",1081=> X"0200",1082=> X"1700",1083=> X"0000",1084=> X"0000",1085=> X"0000",1086=> X"0000",1087=> X"0000",1088=> X"b800",1089=> X"0200",1090=> X"1100",1091=> X"0000",1092=> X"0000",1093=> X"0000",1094=> X"0000",1095=> X"0000",1096=> X"8e00",1097=> X"0200",1098=> X"1100",1099=> X"0000",1100=> X"0000",1101=> X"0000",1102=> X"0000",1103=> X"0000",1104=> X"8380",1105=> X"0200",1106=> X"1100",1107=> X"0000",1108=> X"0000",1109=> X"0000",1110=> X"0000",1111=> X"0000",1112=> X"80e0",1113=> X"0200",1114=> X"1d00",1115=> X"0000",1116=> X"0000",1117=> X"0000",1118=> X"0000",1119=> X"0000",1120=> X"8038",1121=> X"0200",1122=> X"1100",1123=> X"0000",1124=> X"0000",1125=> X"0000",1126=> X"0000",1127=> X"0000",1128=> X"800f",1129=> X"fffc",1130=> X"1100",1131=> X"0000",1132=> X"0000",1133=> X"0000",1134=> X"0000",1135=> X"0000",1136=> X"8000",1137=> X"0004",1138=> X"1100",1139=> X"0000",1140=> X"0000",1141=> X"0000",1142=> X"0000",1143=> X"0000",1144=> X"8000",1145=> X"0004",1146=> X"1700",1147=> X"0000",1148=> X"0000",1149=> X"0000",1150=> X"0000",1151=> X"0000",1152=> X"8000",1153=> X"0004",1154=> X"1100",1155=> X"0000",1156=> X"0000",1157=> X"0000",1158=> X"0000",1159=> X"0000",1160=> X"8000",1161=> X"0004",1162=> X"1100",1163=> X"0000",1164=> X"0000",1165=> X"0000",1166=> X"0000",1167=> X"0000",1168=> X"8000",1169=> X"0004",1170=> X"1100",1171=> X"0000",1172=> X"0000",1173=> X"0000",1174=> X"0000",1175=> X"0000",1176=> X"8000",1177=> X"0004",1178=> X"1d00",1179=> X"0000",1180=> X"0000",1181=> X"0000",1182=> X"0000",1183=> X"0000",1184=> X"8000",1185=> X"0004",1186=> X"0100",1187=> X"0000",1188=> X"0000",1189=> X"0000",1190=> X"0000",1191=> X"0000",1192=> X"ffff",1193=> X"ffff",1194=> X"ff00",1195=> X"0000",1196=> X"0000",1197=> X"0000",1198=> X"0000",1199=> X"0000",1200=> X"0000",1201=> X"0000",1202=> X"0000",1203=> X"0000",1204=> X"0000",1205=> X"0000",1206=> X"0000",1207=> X"0000",1208=> X"0000",1209=> X"0000",1210=> X"0000",1211=> X"0000",1212=> X"0000",1213=> X"0000",1214=> X"0000",1215=> X"0000",1216=> X"0000",1217=> X"0000",1218=> X"0000",1219=> X"0000",1220=> X"0000",1221=> X"0000",1222=> X"0000",1223=> X"0000",1224=> X"0000",1225=> X"0000",1226=> X"0000",1227=> X"0000",1228=> X"0000",1229=> X"0000",1230=> X"0000",1231=> X"0000",1232=> X"0000",1233=> X"0000",1234=> X"0000",1235=> X"0000",1236=> X"0000",1237=> X"0000",1238=> X"0000",1239=> X"0000",1240=> X"0000",1241=> X"0000",1242=> X"0000",1243=> X"0000",1244=> X"0000",1245=> X"0000",1246=> X"0000",1247=> X"0000",1248=> X"0000",1249=> X"0000",1250=> X"0000",1251=> X"0000",1252=> X"0000",1253=> X"0000",1254=> X"0000",1255=> X"0000",1256=> X"0000",1257=> X"0000",1258=> X"0000",1259=> X"0000",1260=> X"0000",1261=> X"0000",1262=> X"0000",1263=> X"0000",1264=> X"0000",1265=> X"0000",1266=> X"0000",1267=> X"0000",1268=> X"0000",1269=> X"0000",1270=> X"0000",1271=> X"0000",1272=> X"0000",1273=> X"0000",1274=> X"0000",1275=> X"0000",1276=> X"0000",1277=> X"0000",1278=> X"0000",1279=> X"0000",
                                        1600=> X"ffff",1601=> X"ffff",1602=> X"ff00",1603=> X"0000",1604=> X"0000",1605=> X"0000",1606=> X"0000",1607=> X"0000",1608=> X"8000",1609=> X"0000",1610=> X"0100",1611=> X"0000",1612=> X"0000",1613=> X"0000",1614=> X"0000",1615=> X"0000",1616=> X"8000",1617=> X"0000",1618=> X"0100",1619=> X"0000",1620=> X"0000",1621=> X"0000",1622=> X"0000",1623=> X"0000",1624=> X"8000",1625=> X"0000",1626=> X"0100",1627=> X"0000",1628=> X"0000",1629=> X"0000",1630=> X"0000",1631=> X"0000",1632=> X"8000",1633=> X"0070",1634=> X"0100",1635=> X"0000",1636=> X"0000",1637=> X"0000",1638=> X"0000",1639=> X"0000",1640=> X"8000",1641=> X"0088",1642=> X"0100",1643=> X"0000",1644=> X"0000",1645=> X"0000",1646=> X"0000",1647=> X"0000",1648=> X"8000",1649=> X"0104",1650=> X"0100",1651=> X"0000",1652=> X"0000",1653=> X"0000",1654=> X"0000",1655=> X"0000",1656=> X"8000",1657=> X"0104",1658=> X"0100",1659=> X"0000",1660=> X"0000",1661=> X"0000",1662=> X"0000",1663=> X"0000",1664=> X"8000",1665=> X"0202",1666=> X"0100",1667=> X"0000",1668=> X"0000",1669=> X"0000",1670=> X"0000",1671=> X"0000",1672=> X"8000",1673=> X"1e02",1674=> X"0100",1675=> X"0000",1676=> X"0000",1677=> X"0000",1678=> X"0000",1679=> X"0000",1680=> X"8000",1681=> X"0202",1682=> X"0100",1683=> X"0000",1684=> X"0000",1685=> X"0000",1686=> X"0000",1687=> X"0000",1688=> X"8000",1689=> X"0202",1690=> X"0100",1691=> X"0000",1692=> X"0000",1693=> X"0000",1694=> X"0000",1695=> X"0000",1696=> X"8000",1697=> X"0202",1698=> X"0100",1699=> X"0000",1700=> X"0000",1701=> X"0000",1702=> X"0000",1703=> X"0000",1704=> X"8fff",1705=> X"fe00",1706=> X"0100",1707=> X"0000",1708=> X"0000",1709=> X"0000",1710=> X"0000",1711=> X"0000",1712=> X"8000",1713=> X"2000",1714=> X"0100",1715=> X"0000",1716=> X"0000",1717=> X"0000",1718=> X"0000",1719=> X"0000",1720=> X"8000",1721=> X"2000",1722=> X"0700",1723=> X"0000",1724=> X"0000",1725=> X"0000",1726=> X"0000",1727=> X"0000",1728=> X"8000",1729=> X"2000",1730=> X"0100",1731=> X"0000",1732=> X"0000",1733=> X"0000",1734=> X"0000",1735=> X"0000",1736=> X"8000",1737=> X"2000",1738=> X"0100",1739=> X"0000",1740=> X"0000",1741=> X"0000",1742=> X"0000",1743=> X"0000",1744=> X"8000",1745=> X"2000",1746=> X"0100",1747=> X"0000",1748=> X"0000",1749=> X"0000",1750=> X"0000",1751=> X"0000",1752=> X"8000",1753=> X"2000",1754=> X"0100",1755=> X"0000",1756=> X"0000",1757=> X"0000",1758=> X"0000",1759=> X"0000",1760=> X"8000",1761=> X"2000",1762=> X"0100",1763=> X"0000",1764=> X"0000",1765=> X"0000",1766=> X"0000",1767=> X"0000",1768=> X"800f",1769=> X"fffc",1770=> X"0100",1771=> X"0000",1772=> X"0000",1773=> X"0000",1774=> X"0000",1775=> X"0000",1776=> X"8038",1777=> X"0000",1778=> X"0100",1779=> X"0000",1780=> X"0000",1781=> X"0000",1782=> X"0000",1783=> X"0000",1784=> X"8068",1785=> X"0000",1786=> X"0700",1787=> X"0000",1788=> X"0000",1789=> X"0000",1790=> X"0000",1791=> X"0000",1792=> X"80c8",1793=> X"0000",1794=> X"0100",1795=> X"0000",1796=> X"0000",1797=> X"0000",1798=> X"0000",1799=> X"0000",1800=> X"8188",1801=> X"0000",1802=> X"0100",1803=> X"0000",1804=> X"0000",1805=> X"0000",1806=> X"0000",1807=> X"0000",1808=> X"8308",1809=> X"0000",1810=> X"0100",1811=> X"0000",1812=> X"0000",1813=> X"0000",1814=> X"0000",1815=> X"0000",1816=> X"8608",1817=> X"0000",1818=> X"0100",1819=> X"0000",1820=> X"0000",1821=> X"0000",1822=> X"0000",1823=> X"0000",1824=> X"8c08",1825=> X"0000",1826=> X"0100",1827=> X"0000",1828=> X"0000",1829=> X"0000",1830=> X"0000",1831=> X"0000",1832=> X"ffff",1833=> X"ffff",1834=> X"ff00",1835=> X"0000",1836=> X"0000",1837=> X"0000",1838=> X"0000",1839=> X"0000",1840=> X"0000",1841=> X"0000",1842=> X"0000",1843=> X"0000",1844=> X"0000",1845=> X"0000",1846=> X"0000",1847=> X"0000",1848=> X"0000",1849=> X"0000",1850=> X"0000",1851=> X"0000",1852=> X"0000",1853=> X"0000",1854=> X"0000",1855=> X"0000",1856=> X"0000",1857=> X"0000",1858=> X"0000",1859=> X"0000",1860=> X"0000",1861=> X"0000",1862=> X"0000",1863=> X"0000",1864=> X"0000",1865=> X"0000",1866=> X"0000",1867=> X"0000",1868=> X"0000",1869=> X"0000",1870=> X"0000",1871=> X"0000",1872=> X"0000",1873=> X"0000",1874=> X"0000",1875=> X"0000",1876=> X"0000",1877=> X"0000",1878=> X"0000",1879=> X"0000",1880=> X"0000",1881=> X"0000",1882=> X"0000",1883=> X"0000",1884=> X"0000",1885=> X"0000",1886=> X"0000",1887=> X"0000",1888=> X"0000",1889=> X"0000",1890=> X"0000",1891=> X"0000",1892=> X"0000",1893=> X"0000",1894=> X"0000",1895=> X"0000",1896=> X"0000",1897=> X"0000",1898=> X"0000",1899=> X"0000",1900=> X"0000",1901=> X"0000",1902=> X"0000",1903=> X"0000",1904=> X"0000",1905=> X"0000",1906=> X"0000",1907=> X"0000",1908=> X"0000",1909=> X"0000",1910=> X"0000",1911=> X"0000",1912=> X"0000",1913=> X"0000",1914=> X"0000",1915=> X"0000",1916=> X"0000",1917=> X"0000",1918=> X"0000",1919=> X"0000",
                                      others=> X"0000");

    -- Micro memory
    type uMem_type is array (0 to 511) of STD_LOGIC_VECTOR(31 downto 0);
    constant uMem : uMem_type := (  0=>X"04100000",
                                    1=>X"03280000",
                                    2=>X"00000400",
                                    3=>X"0A540200",
                                    4=>X"04180000",
                                    5=>X"03500200",
                                    6=>X"04180000",
                                    7=>X"03100000",
                                    8=>X"03500200",
                                    9=>X"05A00600",
                                    10=>X"05100000",
                                    11=>X"0A300600",
                                    12=>X"15000000",
                                    13=>X"4A000000",
                                    14=>X"07A00600",
                                    15=>X"05400600",
                                    16=>X"00002A0F",
                                    17=>X"00000600",
                                    18=>X"0000220F",
                                    19=>X"00000600",
                                    20=>X"0000240F",
                                    21=>X"00000600",
                                    22=>X"00003816",
                                    23=>X"00000600",
                                    24=>X"1A000000",
                                    25=>X"55000600",
                                    26=>X"09100000",
                                    27=>X"04300000",
                                    28=>X"05420600",
                                    29=>X"00010000",
                                    30=>X"09100000",
                                    31=>X"03400600",
                                    32=>X"09100000",
                                    33=>X"0A320600",
                                    34=>X"00010000",
                                    35=>X"09100000",
                                    36=>X"03A00600",
                                    37=>X"05900600",
                                    38=>X"1A000000",
                                    39=>X"55000000",
                                    40=>X"07A00600",
                                    41=>X"05008000",
                                    42=>X"1A00342D",
                                    43=>X"D0004000",
                                    44=>X"0000322B",
                                    45=>X"07A00600",
                                    46=>X"05008000",
                                    47=>X"1A003432",
                                    48=>X"90004000",
                                    49=>X"00003230",
                                    50=>X"07A00600",
                                    51=>X"15000000",
                                    52=>X"6A000000",
                                    53=>X"07A00600",
                                    54=>X"15000000",
                                    55=>X"7A000000",
                                    56=>X"07A00600",
                                    57=>X"04180000",
                                    58=>X"13000000",
                                    59=>X"4A040000",
                                    60=>X"07100000",
                                    61=>X"03500200",
                                    62=>X"0000260F",
                                    63=>X"00000600",
                                    64=>X"0000280F",
                                    65=>X"00000600",
                                    66=>X"30000000",
                                    67=>X"55000000",
                                    68=>X"07A00600",
                                    69=>X"05008000",
                                    70=>X"00003846",
                                    71=>X"00007246",
                                    72=>X"00000600",
                                    511=>X"00003E00",
                                    others=> X"00000000");

    -- uPC
    signal uPC : STD_LOGIC_VECTOR(8 downto 0) := (others=>'0');
    signal SuPC : STD_LOGIC_VECTOR(8 downto 0) := (others=>'0');

    signal ctrlword : STD_LOGIC_VECTOR(31 downto 0) := X"00000000";
    alias cALU : STD_LOGIC_VECTOR(3 downto 0) is ctrlword(31 downto 28);
    alias cTB : STD_LOGIC_VECTOR(3 downto 0) is ctrlword(27 downto 24);
    alias cFB : STD_LOGIC_VECTOR(3 downto 0) is ctrlword(23 downto 20);
    alias cP : STD_LOGIC is ctrlword(19);
    alias cM : STD_LOGIC is ctrlword(18);
    alias cSP : STD_LOGIC_VECTOR(1 downto 0) is ctrlword(17 downto 16);
    alias cLC : STD_LOGIC_VECTOR(1 downto 0) is ctrlword(15 downto 14);
    alias cSEQ : STD_LOGIC_VECTOR(4 downto 0) is ctrlword(13 downto 9);
    alias cADR : STD_LOGIC_VECTOR(8 downto 0) is ctrlword(8 downto 0);

    type K1_type is array (0 to 63) of STD_LOGIC_VECTOR(8 downto 0);
    signal K1 : K1_type := (0=>"000001001", --MOVE
                            1=>"000001010", --STORE
                            2=>"000001100", --ADD
                            3=>"000001111", --BRA
                            4=>"000010000", --BCS
                            5=>"000010010", --BEQ
                            6=>"000010100", --BNE
                            7=>"000010110", --WVS
                            8=>"000011000", --CMP
                            9=>"000011010", --JSR
                            10=>"000011101", --RTS
                            11=>"000100000", --PUSH
                            12=>"000100010", --POP
                            13=>"000100101", --SSP
                            14=>"000100110", --SUB
                            15=>"000101001", --LSR
                            16=>"000101110", --LSL
                            17=>"000110011", --AND
                            18=>"000110110", --OR
                            19=>"000111110", --BMI
                            20=>"001000000", --BPL
                            21=>"001000010", --INV
                            22=>"001000101", --LWVS  
                            others=>"111111111"); --HULT

    type K2_type is array (0 to 3) of STD_LOGIC_VECTOR(8 downto 0);
    signal K2 : K2_type := (0=>"000000011", --reg-reg
                            1=>"000000100", --imm
                            2=>"000000110", --indir
                            3=>"000111001", --index
                            others=>"000000000");

    type gr_array is array (0 to 15) of STD_LOGIC_VECTOR(15 downto 0);
    signal rGR : gr_array := (others=> X"0000");

    signal tempGR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal tempPM : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal tempMM : STD_LOGIC_VECTOR(15 downto 0) := X"0000";


    ---------- DEBUG --------
    signal old_step : STD_LOGIC := '0';

begin
    ctrlword <= uMem(conv_integer(uPC));

    led_driver: leddriver port map (clk, rst, seg, an, led, rGR(2), rGR(5)(0) & rGR(4)(0) & "00000" & rGR(3)(0)); --rGR(2) 7-seg, rGR(3) leds
    --led_driver: leddriver port map (clk, rst, seg, an, led, rGR(2), rGR(5)(7 downto 0)); --rGR(2) 7-seg, rGR(3) leds
    alu_instance: alu port map(clk, cALU, rAR, databus, rAR, fC, fZ, fN, fO);
    

    -- *****************************
    -- * CONTROL UNIT              *
    -- *****************************
    process(clk) begin
        if rising_edge(clk) then
            
            -- rst
            if rst = '1' then
                rPC <= X"0000";
                uPC <= "000000000";
            else

                -- LC control
                case cLC is
                    when "01" => rLC <= rLC - 1;
                    when "10" => rLC <= databus(7 downto 0);
                    when "11" => rLC <= cADR(7 downto 0);
                    when others => null;
                end case;

                -- P control
                if cP = '1' then
                    rPC <= rPC + 1; 
                end if;

                -- SP control
                case cSP is
                    when "01" => rSP <= rSP + 1;
                    when "10" => rSP <= rSP - 1;
                    when others => null;
                end case;

                -- SEQ
                case cSEQ is
                    when "00000" => uPC <= uPC + 1;
                    when "00001" => uPC <= K1(conv_integer(rIR(15 downto 10)));
                    when "00010" => uPC <= K2(conv_integer(rIR(9 downto 8)));
                    when "00011" => uPC <= "000000000";
                    when "10000" => uPC <= cADR;
                    when "10001" => if fZ = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10010" => if fZ = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10011" => if fN = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10100" => if fN = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10101" => if fC = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10110" => if fC = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10111" => if fO = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11000" => if fO = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11001" => if fL = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11010" => if fL = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11011" => if fV = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11100" => if fV = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11101" => 
                        uPC <= cADR; 
                        SuPC <= uPC+1;
                    when "11110" => uPC <= SuPC;
                    when "11111" => null;
                    when others => null;
                end case;
                
                -- FROM BUS
                case cFB is
                    when "0001" => rASR <= databus;
                    when "0010" => rIR <= databus;
                    when "0011" => 
                        if (rASR(15) = '0') then
                            PrimMem(conv_integer(rASR)) <= databus;
                        elsif (rASR(15 downto 12) = X"9") then -- VR
                            vr_i <= databus;
                        end if;
                    when "0100" => rPC <= databus;
                    when "0101" => rDR <= databus;
                    when "0110" => null; -- can't write to uM
                    when "0111" => null; -- can't write to AR
                    when "1000" => rHR <= databus;
                    when "1001" => rSP <= databus;
                    when "1010" => 
                        if cM = '0' then 
                            rGR(conv_integer(rIR(7 downto 4))) <= databus;
                        else
                            rGR(conv_integer(rIR(3 downto 0))) <= databus;
                        end if;
                    when others => null;
                end case;
            end if;
        end if;
    end process;

    with rLC select
    fL <= '0' when X"00",
          '1' when others;

    --process(cFB, rASR, databus) begin
    process(clk) begin
        if rising_edge(clk) then
            if cFB = "0011" and rASR(15 downto 12) = X"9" then -- 9xxx address
                vr_we <= '1';
                --vr_i <= databus;
            else
                vr_we <= '0';
            end if;
        end if;
    end process;

    vr_addr <= rASR(4 downto 0);

    -- TO BUS
    with cTB select
    databus <= rASR when "0001",
                rIR when "0010",
                tempPM when "0011", -- PM/MM
                rPC when "0100",
                rDR when "0101",
                --uMem(conv_integer(uPC)) when "0110",
                rAR when "0111",
                rHR when "1000",
                rSP when "1001",
                tempGR when "1010",
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                --vr_o when "1011",
                X"0000" when others;

    -- PM/MemMap
    with rASR(15) select
    tempPM <= PrimMem(conv_integer(rASR)) when '0',
              tempMM when others;

    -- MemMap
    with rASR select
    tempMM <= "000000000000000" & up when X"8000",
              "000000000000000" & right when X"8001",
              "000000000000000" & down when X"8002",
              "000000000000000" & left when X"8003",
              X"00" & sw when X"8004",
              --X"00" & ledval when X"A000",
              --value when X"A001",
              vr_o when X"9000",vr_o when X"9001",vr_o when X"9002",vr_o when X"9003",
              vr_o when X"9004",vr_o when X"9005",vr_o when X"9006",vr_o when X"9007",
              vr_o when X"9008",vr_o when X"9009",vr_o when X"900A",vr_o when X"900B",
              vr_o when X"900C",vr_o when X"900D",vr_o when X"900E",vr_o when X"900F",
              vr_o when X"9010",vr_o when X"9011",vr_o when X"9012",vr_o when X"9013",
              vr_o when X"9014",vr_o when X"9015",vr_o when X"9016",vr_o when X"9017",
              vr_o when X"9018",vr_o when X"9019",vr_o when X"901A",vr_o when X"901B",
              vr_o when X"901C",vr_o when X"901D",vr_o when X"901E",vr_o when X"901F",
              X"EEEE" when others;

    -- M bit
    with cM select
    tempGR <= rGR(conv_integer(rIR(7 downto 4))) when '0',
              rGR(conv_integer(rIR(3 downto 0))) when others;

end cpu_one;
