library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity alu is
    Port (  clk : in STD_LOGIC;
            op : in STD_LOGIC_VECTOR(3 downto 0);
            A, B : in STD_LOGIC_VECTOR(15 downto 0);
            result : out STD_LOGIC_VECTOR(15 downto 0);
            carry, zero, negative, overflow : out STD_LOGIC);
end alu;

architecture alu_one of alu is
    signal value : STD_LOGIC_VECTOR(16 downto 0) := "00000000000000000";
    signal useflag : STD_LOGIC := '0';

begin
    process(A, B, op) begin
        case op is
            when "0001" => value <= '0' & B; --databus
                           useflag <= '1';
            when "0011" => value <= "00000000000000000"; --nollställ
                           useflag <= '1';
            when "0100" => value <= STD_LOGIC_VECTOR('0' & unsigned(A) + unsigned(B)); --add
                           useflag <= '1';
            when "0101" => value <= ('0' & A) - B; --sub
                           useflag <= '1';
            when "0110" => value <= '0' & A and '0' & B; -- and
                           useflag <= '1';
            when "0111" => value <= '0' & A or '0' & B; -- or
                           useflag <= '1';
            when "1000" => value <= STD_LOGIC_VECTOR('0' & unsigned(A) + unsigned(B)); --add noflag
                           useflag <= '0';
            when "1001" => value <= a & '0'; -- ASL/LSL
                           useflag <= '1';
            when "1011" => value <= a(0) & a(15) & a(15 downto 1); -- ASR
                           useflag <= '1';
            when "1101" => value <= a(0) & '0' & a(15 downto 1); -- LSR
                           useflag <= '1';
            when others => value <= '0' & A; -- AR
                           useflag <= '0';
        end case;
    end process;
    
    process(clk) begin
    --process(value, useflag) begin
        if rising_edge(clk) then
            result <= value(15 downto 0);
            if useflag = '1' then
                if value(15 downto 0) = X"0000" then
                    zero <= '1';
                else
                    zero <= '0';
                end if;
                if value(16) = '1' then carry <= '1';
                else carry <= '0'; 
                end if;
                if value(15) = '1' then negative <= '1'; 
                else negative <= '0'; 
                end if;
                if value(16) /= value(15) then overflow <= '1';
                else overflow <= '0';
                end if;
            end if; 
        end if;
    end process;
end alu_one;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity cpu is
    Port (clk,rst : in  STD_LOGIC;
        sw: in STD_LOGIC_VECTOR(7 downto 0);
        seg: out  STD_LOGIC_VECTOR(7 downto 0);
        an : out  STD_LOGIC_VECTOR (3 downto 0);
        led : out STD_LOGIC_VECTOR (7 downto 0);
        vr_we : out STD_LOGIC;
        vr_addr : out STD_LOGIC_VECTOR(4 downto 0);
        vr_i : out STD_LOGIC_VECTOR(15 downto 0);
        vr_o : in STD_LOGIC_VECTOR(15 downto 0);
        fV: in STD_LOGIC;
        up, right, down, left : in STD_LOGIC);
end cpu;

architecture cpu_one of cpu is

    component leddriver
        Port ( clk,rst : in  STD_LOGIC;
           seg : out  STD_LOGIC_VECTOR(7 downto 0);
           an : out  STD_LOGIC_VECTOR (3 downto 0);
           led : out STD_LOGIC_VECTOR (7 downto 0);
           value : in  STD_LOGIC_VECTOR (15 downto 0);
           ledval : in STD_LOGIC_VECTOR (7 downto 0));
    end component;

    component alu
        Port (clk : in STD_LOGIC;
            op : in STD_LOGIC_VECTOR(3 downto 0);
            A, B : in STD_LOGIC_VECTOR(15 downto 0);
            result : out STD_LOGIC_VECTOR(15 downto 0);
            carry, zero, negative, overflow : out STD_LOGIC);
    end component;

    signal databus : STD_LOGIC_VECTOR(15 downto 0) := X"0000";

    -- Registers
    signal rASR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rIR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rPC : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rDR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rAR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rHR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rSP : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rLC : STD_LOGIC_VECTOR(7 downto 0) := X"00";

    -- Flags
    signal fZ : STD_LOGIC := '1';
    signal fN : STD_LOGIC := '0';
    signal fC : STD_LOGIC := '0';
    signal fO : STD_LOGIC := '0';
    signal fL : STD_LOGIC := '0';

    -- Primary memory
    type PrimMem_type is array (0 to 2047) of STD_LOGIC_VECTOR(15 downto 0);
    signal PrimMem : PrimMem_type := (  0=> X"0100",1=> X"0000",2=> X"0110",3=> X"00d0",4=> X"0140",5=> X"00f0",6=> X"0120",7=> X"0001",8=> X"0130",9=> X"0002",10=> X"0540",11=> X"0022",12=> X"0510",13=> X"0023",14=> X"0500",15=> X"0024",16=> X"0500",17=> X"0025",18=> X"0500",19=> X"0026",20=> X"0500",21=> X"0027",22=> X"0500",23=> X"0028",24=> X"0500",25=> X"002d",26=> X"0500",27=> X"002e",28=> X"0520",29=> X"002f",30=> X"0530",31=> X"0030",32=> X"0d00",33=> X"004a",34=> X"0000",35=> X"0000",36=> X"0000",37=> X"0000",38=> X"0000",39=> X"0000",40=> X"0000",41=> X"0000",42=> X"0000",43=> X"0000",44=> X"0000",45=> X"0000",46=> X"0000",47=> X"0000",48=> X"0000",49=> X"0000",50=> X"0000",51=> X"0000",52=> X"0000",53=> X"0000",54=> X"0002",55=> X"0000",56=> X"0000",57=> X"0000",58=> X"fffc",59=> X"0000",60=> X"0000",61=> X"0000",62=> X"0000",63=> X"0000",64=> X"00e0",65=> X"01a0",66=> X"01f0",67=> X"0140",68=> X"00c0",69=> X"00c0",70=> X"0130",71=> X"01c0",72=> X"0640",73=> X"0500",74=> X"3500",75=> X"07ff",76=> X"2500",77=> X"0073",78=> X"2500",79=> X"0080",80=> X"2500",81=> X"00d5",82=> X"2500",83=> X"010c",84=> X"2500",85=> X"0149",86=> X"2500",87=> X"0168",88=> X"0200",89=> X"0022",90=> X"4500",91=> X"0fff",92=> X"0500",93=> X"0022",94=> X"2500",95=> X"0187",96=> X"2500",97=> X"01f4",98=> X"2500",99=> X"0325",100=> X"2500",101=> X"036a",102=> X"2500",103=> X"037d",104=> X"0220",105=> X"003e",106=> X"0230",107=> X"0022",108=> X"0240",109=> X"002d",110=> X"0250",111=> X"0025",112=> X"1c00",113=> X"0d00",114=> X"004c",115=> X"2d00",116=> X"0000",117=> X"0200",118=> X"003d",119=> X"0900",120=> X"0001",121=> X"4500",122=> X"0003",123=> X"0500",124=> X"003d",125=> X"3100",126=> X"0000",127=> X"2800",128=> X"2d00",129=> X"0000",130=> X"2d10",131=> X"0000",132=> X"0200",133=> X"8004",134=> X"4500",135=> X"0001",136=> X"0500",137=> X"0024",138=> X"0200",139=> X"8000",140=> X"0210",141=> X"0033",142=> X"4a10",143=> X"0034",144=> X"0801",145=> X"2100",146=> X"0002",147=> X"1900",148=> X"009d",149=> X"0100",150=> X"0020",151=> X"0500",152=> X"0028",153=> X"0100",154=> X"0000",155=> X"0500",156=> X"0027",157=> X"0200",158=> X"8001",159=> X"0210",160=> X"8003",161=> X"2001",162=> X"4d00",163=> X"00b0",164=> X"1500",165=> X"00ba",166=> X"0110",167=> X"0002",168=> X"0510",169=> X"002e",170=> X"0110",171=> X"0001",172=> X"0510",173=> X"002d",174=> X"0d00",175=> X"00d0",176=> X"0110",177=> X"0002",178=> X"0510",179=> X"002e",180=> X"0110",181=> X"0000",182=> X"0510",183=> X"002d",184=> X"0d00",185=> X"00d0",186=> X"0210",187=> X"0026",188=> X"2110",189=> X"0000",190=> X"1500",191=> X"00cc",192=> X"5610",193=> X"0025",194=> X"0910",195=> X"0001",196=> X"0510",197=> X"002d",198=> X"0110",199=> X"0001",200=> X"0510",201=> X"002e",202=> X"0d00",203=> X"00d0",204=> X"0110",205=> X"0000",206=> X"0510",207=> X"002e",208=> X"3110",209=> X"0000",210=> X"3100",211=> X"0000",212=> X"2800",213=> X"2d00",214=> X"0000",215=> X"2d10",216=> X"0000",217=> X"0200",218=> X"0025",219=> X"2200",220=> X"002d",221=> X"1500",222=> X"00e1",223=> X"1900",224=> X"00e9",225=> X"0200",226=> X"0026",227=> X"0a00",228=> X"002e",229=> X"0500",230=> X"0026",231=> X"0d00",232=> X"00fd",233=> X"0200",234=> X"0026",235=> X"3a00",236=> X"002e",237=> X"4d00",238=> X"00f3",239=> X"0500",240=> X"0026",241=> X"0d00",242=> X"00fd",243=> X"5600",244=> X"0026",245=> X"0500",246=> X"0026",247=> X"5600",248=> X"0025",249=> X"0900",250=> X"0001",251=> X"0500",252=> X"0025",253=> X"0200",254=> X"0026",255=> X"2100",256=> X"0018",257=> X"4d00",258=> X"0107",259=> X"0100",260=> X"0018",261=> X"0500",262=> X"0026",263=> X"3110",264=> X"0000",265=> X"3100",266=> X"0000",267=> X"2800",268=> X"2d00",269=> X"0000",270=> X"2d10",271=> X"0000",272=> X"0200",273=> X"0027",274=> X"2200",275=> X"002f",276=> X"1500",277=> X"0118",278=> X"1900",279=> X"0120",280=> X"0200",281=> X"0028",282=> X"0a00",283=> X"0030",284=> X"0500",285=> X"0028",286=> X"0d00",287=> X"0134",288=> X"0200",289=> X"0028",290=> X"3a00",291=> X"0030",292=> X"4d00",293=> X"012a",294=> X"0500",295=> X"0028",296=> X"0d00",297=> X"0134",298=> X"5600",299=> X"0028",300=> X"0500",301=> X"0028",302=> X"5600",303=> X"0027",304=> X"0900",305=> X"0001",306=> X"0500",307=> X"0027",308=> X"0200",309=> X"0027",310=> X"2100",311=> X"0001",312=> X"1900",313=> X"0144",314=> X"0200",315=> X"0028",316=> X"2100",317=> X"0020",318=> X"4d00",319=> X"0144",320=> X"0100",321=> X"0020",322=> X"0500",323=> X"0028",324=> X"3110",325=> X"0000",326=> X"3100",327=> X"0000",328=> X"2800",329=> X"2d00",330=> X"0000",331=> X"2d10",332=> X"0000",333=> X"2d80",334=> X"0000",335=> X"0200",336=> X"0026",337=> X"0210",338=> X"0022",339=> X"3d00",340=> X"0003",341=> X"0280",342=> X"0025",343=> X"2180",344=> X"0001",345=> X"1900",346=> X"015e",347=> X"0810",348=> X"0d00",349=> X"015f",350=> X"3810",351=> X"0510",352=> X"0022",353=> X"3180",354=> X"0000",355=> X"3110",356=> X"0000",357=> X"3100",358=> X"0000",359=> X"2800",360=> X"2d00",361=> X"0000",362=> X"2d10",363=> X"0000",364=> X"2d80",365=> X"0000",366=> X"0200",367=> X"0028",368=> X"0210",369=> X"0023",370=> X"3d00",371=> X"0003",372=> X"0280",373=> X"0027",374=> X"2180",375=> X"0001",376=> X"1900",377=> X"017d",378=> X"0810",379=> X"0d00",380=> X"017e",381=> X"3810",382=> X"0510",383=> X"0023",384=> X"3180",385=> X"0000",386=> X"3110",387=> X"0000",388=> X"3100",389=> X"0000",390=> X"2800",391=> X"2d00",392=> X"0000",393=> X"2d10",394=> X"0000",395=> X"2d20",396=> X"0000",397=> X"0200",398=> X"0022",399=> X"0210",400=> X"0023",401=> X"2500",402=> X"01bc",403=> X"0500",404=> X"0031",405=> X"0200",406=> X"0022",407=> X"0900",408=> X"000f",409=> X"0210",410=> X"0023",411=> X"2500",412=> X"01bc",413=> X"0500",414=> X"0032",415=> X"0200",416=> X"0022",417=> X"0210",418=> X"0023",419=> X"0910",420=> X"000f",421=> X"2500",422=> X"01bc",423=> X"0500",424=> X"0033",425=> X"0200",426=> X"0022",427=> X"0900",428=> X"000f",429=> X"0210",430=> X"0023",431=> X"0910",432=> X"000f",433=> X"2500",434=> X"01bc",435=> X"0500",436=> X"0034",437=> X"3120",438=> X"0000",439=> X"3110",440=> X"0000",441=> X"3100",442=> X"0000",443=> X"2800",444=> X"2d20",445=> X"0000",446=> X"2d30",447=> X"0000",448=> X"2d40",449=> X"0000",450=> X"2df0",451=> X"0000",452=> X"3d00",453=> X"0004",454=> X"3d10",455=> X"0004",456=> X"0050",457=> X"3d00",458=> X"0004",459=> X"4500",460=> X"0007",461=> X"4110",462=> X"0003",463=> X"0801",464=> X"02f0",465=> X"0024",466=> X"03ff",467=> X"0048",468=> X"08f0",469=> X"032f",470=> X"0000",471=> X"0005",472=> X"4500",473=> X"000f",474=> X"0130",475=> X"000f",476=> X"3830",477=> X"0140",478=> X"0001",479=> X"4043",480=> X"4424",481=> X"2120",482=> X"0000",483=> X"1500",484=> X"01e9",485=> X"0100",486=> X"0001",487=> X"0d00",488=> X"01eb",489=> X"0100",490=> X"0000",491=> X"31f0",492=> X"0000",493=> X"3140",494=> X"0000",495=> X"3130",496=> X"0000",497=> X"3120",498=> X"0000",499=> X"2800",500=> X"2d00",501=> X"0000",502=> X"2d10",503=> X"0000",504=> X"2d20",505=> X"0000",506=> X"0200",507=> X"0031",508=> X"2100",509=> X"0001",510=> X"1500",511=> X"0214",512=> X"0200",513=> X"0032",514=> X"2100",515=> X"0001",516=> X"1500",517=> X"0222",518=> X"0200",519=> X"0033",520=> X"2100",521=> X"0001",522=> X"1500",523=> X"022a",524=> X"0200",525=> X"0034",526=> X"2100",527=> X"0001",528=> X"1500",529=> X"031a",530=> X"0d00",531=> X"031e",532=> X"0200",533=> X"0032",534=> X"2100",535=> X"0001",536=> X"1500",537=> X"0232",538=> X"0200",539=> X"0033",540=> X"2100",541=> X"0001",542=> X"1500",543=> X"0250",544=> X"0d00",545=> X"02f8",546=> X"0200",547=> X"0034",548=> X"2100",549=> X"0001",550=> X"1500",551=> X"0268",552=> X"0d00",553=> X"030a",554=> X"0200",555=> X"0034",556=> X"2100",557=> X"0001",558=> X"1500",559=> X"027d",560=> X"0d00",561=> X"0318",562=> X"0100",563=> X"0000",564=> X"0600",565=> X"0028",566=> X"0200",567=> X"0033",568=> X"2100",569=> X"0001",570=> X"1500",571=> X"028c",572=> X"0200",573=> X"0034",574=> X"2100",575=> X"0001",576=> X"1500",577=> X"02aa",578=> X"0210",579=> X"0023",580=> X"4510",581=> X"000f",582=> X"0220",583=> X"0023",584=> X"0130",585=> X"0010",586=> X"3831",587=> X"0823",588=> X"0520",589=> X"0023",590=> X"0d00",591=> X"031e",592=> X"0100",593=> X"0000",594=> X"0600",595=> X"0026",596=> X"0200",597=> X"0034",598=> X"2100",599=> X"0001",600=> X"1500",601=> X"02c5",602=> X"0210",603=> X"0022",604=> X"4510",605=> X"000f",606=> X"0220",607=> X"0022",608=> X"0130",609=> X"0010",610=> X"3831",611=> X"0823",612=> X"0520",613=> X"0022",614=> X"0d00",615=> X"031e",616=> X"0100",617=> X"0000",618=> X"0600",619=> X"0026",620=> X"0200",621=> X"0033",622=> X"2100",623=> X"0001",624=> X"1500",625=> X"02e0",626=> X"0210",627=> X"0022",628=> X"4510",629=> X"000f",630=> X"0220",631=> X"0022",632=> X"3821",633=> X"0520",634=> X"0022",635=> X"0d00",636=> X"031e",637=> X"0100",638=> X"0000",639=> X"0600",640=> X"0028",641=> X"0210",642=> X"0023",643=> X"4510",644=> X"000f",645=> X"0220",646=> X"0023",647=> X"3821",648=> X"0520",649=> X"0023",650=> X"0d00",651=> X"031e",652=> X"0210",653=> X"0023",654=> X"4510",655=> X"000f",656=> X"0220",657=> X"0023",658=> X"0130",659=> X"0010",660=> X"3831",661=> X"0823",662=> X"0520",663=> X"0023",664=> X"0100",665=> X"0000",666=> X"0600",667=> X"0026",668=> X"0210",669=> X"0022",670=> X"4510",671=> X"000f",672=> X"0220",673=> X"0022",674=> X"0130",675=> X"0010",676=> X"3831",677=> X"0823",678=> X"0520",679=> X"0022",680=> X"0d00",681=> X"031e",682=> X"0210",683=> X"0023",684=> X"4510",685=> X"000f",686=> X"0220",687=> X"0023",688=> X"0130",689=> X"0010",690=> X"3831",691=> X"0823",692=> X"0520",693=> X"0023",694=> X"0100",695=> X"0000",696=> X"0600",697=> X"0026",698=> X"0210",699=> X"0022",700=> X"4510",701=> X"000f",702=> X"0220",703=> X"0022",704=> X"3821",705=> X"0520",706=> X"0022",707=> X"0d00",708=> X"031e",709=> X"0210",710=> X"0022",711=> X"4510",712=> X"000f",713=> X"0220",714=> X"0022",715=> X"0130",716=> X"0010",717=> X"3831",718=> X"0823",719=> X"0520",720=> X"0022",721=> X"0100",722=> X"0000",723=> X"0600",724=> X"0028",725=> X"0210",726=> X"0023",727=> X"4510",728=> X"000f",729=> X"0220",730=> X"0023",731=> X"3821",732=> X"0520",733=> X"0023",734=> X"0d00",735=> X"031e",736=> X"0210",737=> X"0022",738=> X"4510",739=> X"000f",740=> X"0220",741=> X"0022",742=> X"3821",743=> X"0520",744=> X"0022",745=> X"0100",746=> X"0000",747=> X"0600",748=> X"0028",749=> X"0210",750=> X"0023",751=> X"4510",752=> X"000f",753=> X"0220",754=> X"0023",755=> X"3821",756=> X"0520",757=> X"0023",758=> X"0d00",759=> X"031e",760=> X"0100",761=> X"0000",762=> X"0600",763=> X"0028",764=> X"0210",765=> X"0023",766=> X"4510",767=> X"000f",768=> X"0220",769=> X"0023",770=> X"0130",771=> X"0010",772=> X"3831",773=> X"0823",774=> X"0520",775=> X"0023",776=> X"0d00",777=> X"031e",778=> X"0210",779=> X"0023",780=> X"4510",781=> X"000f",782=> X"0220",783=> X"0023",784=> X"0130",785=> X"0010",786=> X"3831",787=> X"0823",788=> X"0520",789=> X"0023",790=> X"0d00",791=> X"031e",792=> X"0d00",793=> X"027d",794=> X"0d00",795=> X"027d",796=> X"0d00",797=> X"031e",798=> X"3120",799=> X"0000",800=> X"3110",801=> X"0000",802=> X"3100",803=> X"0000",804=> X"2800",805=> X"2d00",806=> X"0000",807=> X"2d10",808=> X"0000",809=> X"2df0",810=> X"0000",811=> X"02f0",812=> X"003f",813=> X"030f",814=> X"0040",815=> X"3d00",816=> X"0004",817=> X"0210",818=> X"0022",819=> X"3d10",820=> X"0004",821=> X"2001",822=> X"1500",823=> X"033f",824=> X"0910",825=> X"0001",826=> X"2001",827=> X"1500",828=> X"033f",829=> X"0d00",830=> X"0363",831=> X"030f",832=> X"0044",833=> X"3d00",834=> X"0004",835=> X"0210",836=> X"0023",837=> X"3d10",838=> X"0004",839=> X"2001",840=> X"1500",841=> X"0351",842=> X"0910",843=> X"0001",844=> X"2001",845=> X"1500",846=> X"0351",847=> X"0d00",848=> X"0363",849=> X"0200",850=> X"003e",851=> X"0900",852=> X"0001",853=> X"0500",854=> X"003e",855=> X"0200",856=> X"003d",857=> X"2200",858=> X"003f",859=> X"1900",860=> X"0361",861=> X"0900",862=> X"0001",863=> X"4500",864=> X"0003",865=> X"0500",866=> X"003f",867=> X"31f0",868=> X"0000",869=> X"3110",870=> X"0000",871=> X"3100",872=> X"0000",873=> X"2800",874=> X"2d00",875=> X"0000",876=> X"0200",877=> X"0022",878=> X"3d00",879=> X"0003",880=> X"5400",881=> X"0500",882=> X"0037",883=> X"0200",884=> X"0022",885=> X"3d00",886=> X"0004",887=> X"5400",888=> X"0500",889=> X"0038",890=> X"3100",891=> X"0000",892=> X"2800",893=> X"2d00",894=> X"0000",895=> X"2df0",896=> X"0000",897=> X"02f0",898=> X"0024",899=> X"0200",900=> X"0022",901=> X"0b0f",902=> X"0035",903=> X"0500",904=> X"9000",905=> X"0200",906=> X"0023",907=> X"0b0f",908=> X"0039",909=> X"0500",910=> X"9001",911=> X"0200",912=> X"0024",913=> X"4100",914=> X"000e",915=> X"0500",916=> X"901a",917=> X"0200",918=> X"0035",919=> X"0500",920=> X"9010",921=> X"0200",922=> X"0039",923=> X"0500",924=> X"9011",925=> X"0200",926=> X"0036",927=> X"0500",928=> X"9012",929=> X"0200",930=> X"003a",931=> X"0500",932=> X"9013",933=> X"0200",934=> X"0037",935=> X"0500",936=> X"9014",937=> X"0200",938=> X"003b",939=> X"0500",940=> X"9015",941=> X"0200",942=> X"0038",943=> X"0500",944=> X"9016",945=> X"0200",946=> X"003c",947=> X"0500",948=> X"9017",949=> X"02f0",950=> X"003f",951=> X"030f",952=> X"0040",953=> X"0500",954=> X"9002",955=> X"030f",956=> X"0044",957=> X"0500",958=> X"9003",959=> X"0100",960=> X"0001",961=> X"4100",962=> X"0008",963=> X"0500",964=> X"9018",965=> X"31f0",966=> X"0000",967=> X"3100",968=> X"0000",969=> X"2800",970=> X"2d00",971=> X"0000",972=> X"0200",973=> X"0023",974=> X"3a00",975=> X"8000",976=> X"0a00",977=> X"8002",978=> X"0500",979=> X"0023",980=> X"0200",981=> X"0022",982=> X"0a00",983=> X"8001",984=> X"3a00",985=> X"8003",986=> X"0500",987=> X"0022",988=> X"3100",989=> X"0000",990=> X"2800",
                                        1280=> X"ffff",1281=> X"ffff",1282=> X"ff00",1283=> X"0000",1284=> X"0000",1285=> X"0000",1286=> X"0000",1287=> X"0000",1288=> X"8000",1289=> X"0000",1290=> X"0100",1291=> X"0000",1292=> X"0000",1293=> X"0000",1294=> X"0000",1295=> X"0000",1296=> X"8000",1297=> X"0000",1298=> X"0100",1299=> X"0000",1300=> X"0000",1301=> X"0000",1302=> X"0000",1303=> X"0000",1304=> X"8000",1305=> X"0000",1306=> X"0100",1307=> X"0000",1308=> X"0000",1309=> X"0000",1310=> X"0000",1311=> X"0000",1312=> X"800f",1313=> X"8000",1314=> X"0100",1315=> X"0000",1316=> X"0000",1317=> X"0000",1318=> X"0000",1319=> X"0000",1320=> X"8018",1321=> X"c000",1322=> X"0100",1323=> X"0000",1324=> X"0000",1325=> X"0000",1326=> X"0000",1327=> X"0000",1328=> X"8010",1329=> X"4000",1330=> X"0100",1331=> X"0000",1332=> X"0000",1333=> X"0000",1334=> X"0000",1335=> X"0000",1336=> X"8030",1337=> X"6000",1338=> X"0100",1339=> X"0000",1340=> X"0000",1341=> X"0000",1342=> X"0000",1343=> X"0000",1344=> X"8020",1345=> X"2000",1346=> X"0100",1347=> X"0000",1348=> X"0000",1349=> X"0000",1350=> X"0000",1351=> X"0000",1352=> X"8020",1353=> X"3c00",1354=> X"0100",1355=> X"0000",1356=> X"0000",1357=> X"0000",1358=> X"0000",1359=> X"0000",1360=> X"8020",1361=> X"2000",1362=> X"0100",1363=> X"0000",1364=> X"0000",1365=> X"0000",1366=> X"0000",1367=> X"0000",1368=> X"8020",1369=> X"2000",1370=> X"1d00",1371=> X"0000",1372=> X"0000",1373=> X"0000",1374=> X"0000",1375=> X"0000",1376=> X"8020",1377=> X"2000",1378=> X"1100",1379=> X"0000",1380=> X"0000",1381=> X"0000",1382=> X"0000",1383=> X"0000",1384=> X"8000",1385=> X"03ff",1386=> X"f100",1387=> X"0000",1388=> X"0000",1389=> X"0000",1390=> X"0000",1391=> X"0000",1392=> X"8000",1393=> X"0200",1394=> X"1100",1395=> X"0000",1396=> X"0000",1397=> X"0000",1398=> X"0000",1399=> X"0000",1400=> X"e000",1401=> X"0200",1402=> X"1700",1403=> X"0000",1404=> X"0000",1405=> X"0000",1406=> X"0000",1407=> X"0000",1408=> X"b800",1409=> X"0200",1410=> X"1100",1411=> X"0000",1412=> X"0000",1413=> X"0000",1414=> X"0000",1415=> X"0000",1416=> X"8e00",1417=> X"0200",1418=> X"1100",1419=> X"0000",1420=> X"0000",1421=> X"0000",1422=> X"0000",1423=> X"0000",1424=> X"8380",1425=> X"0200",1426=> X"1100",1427=> X"0000",1428=> X"0000",1429=> X"0000",1430=> X"0000",1431=> X"0000",1432=> X"80e0",1433=> X"0200",1434=> X"1d00",1435=> X"0000",1436=> X"0000",1437=> X"0000",1438=> X"0000",1439=> X"0000",1440=> X"8038",1441=> X"0200",1442=> X"1100",1443=> X"0000",1444=> X"0000",1445=> X"0000",1446=> X"0000",1447=> X"0000",1448=> X"800f",1449=> X"fffc",1450=> X"1100",1451=> X"0000",1452=> X"0000",1453=> X"0000",1454=> X"0000",1455=> X"0000",1456=> X"8000",1457=> X"0004",1458=> X"1100",1459=> X"0000",1460=> X"0000",1461=> X"0000",1462=> X"0000",1463=> X"0000",1464=> X"8000",1465=> X"0004",1466=> X"1700",1467=> X"0000",1468=> X"0000",1469=> X"0000",1470=> X"0000",1471=> X"0000",1472=> X"8000",1473=> X"0004",1474=> X"1100",1475=> X"0000",1476=> X"0000",1477=> X"0000",1478=> X"0000",1479=> X"0000",1480=> X"8000",1481=> X"0004",1482=> X"1100",1483=> X"0000",1484=> X"0000",1485=> X"0000",1486=> X"0000",1487=> X"0000",1488=> X"8000",1489=> X"0004",1490=> X"1100",1491=> X"0000",1492=> X"0000",1493=> X"0000",1494=> X"0000",1495=> X"0000",1496=> X"8000",1497=> X"0004",1498=> X"1d00",1499=> X"0000",1500=> X"0000",1501=> X"0000",1502=> X"0000",1503=> X"0000",1504=> X"8000",1505=> X"0004",1506=> X"0100",1507=> X"0000",1508=> X"0000",1509=> X"0000",1510=> X"0000",1511=> X"0000",1512=> X"ffff",1513=> X"ffff",1514=> X"ff00",1515=> X"0000",1516=> X"0000",1517=> X"0000",1518=> X"0000",1519=> X"0000",1520=> X"0000",1521=> X"0000",1522=> X"0000",1523=> X"0000",1524=> X"0000",1525=> X"0000",1526=> X"0000",1527=> X"0000",1528=> X"0000",1529=> X"0000",1530=> X"0000",1531=> X"0000",1532=> X"0000",1533=> X"0000",1534=> X"0000",1535=> X"0000",1536=> X"0000",1537=> X"0000",1538=> X"0000",1539=> X"0000",1540=> X"0000",1541=> X"0000",1542=> X"0000",1543=> X"0000",1544=> X"0000",1545=> X"0000",1546=> X"0000",1547=> X"0000",1548=> X"0000",1549=> X"0000",1550=> X"0000",1551=> X"0000",1552=> X"0000",1553=> X"0000",1554=> X"0000",1555=> X"0000",1556=> X"0000",1557=> X"0000",1558=> X"0000",1559=> X"0000",1560=> X"0000",1561=> X"0000",1562=> X"0000",1563=> X"0000",1564=> X"0000",1565=> X"0000",1566=> X"0000",1567=> X"0000",1568=> X"0000",1569=> X"0000",1570=> X"0000",1571=> X"0000",1572=> X"0000",1573=> X"0000",1574=> X"0000",1575=> X"0000",1576=> X"0000",1577=> X"0000",1578=> X"0000",1579=> X"0000",1580=> X"0000",1581=> X"0000",1582=> X"0000",1583=> X"0000",1584=> X"0000",1585=> X"0000",1586=> X"0000",1587=> X"0000",1588=> X"0000",1589=> X"0000",1590=> X"0000",1591=> X"0000",1592=> X"0000",1593=> X"0000",1594=> X"0000",1595=> X"0000",1596=> X"0000",1597=> X"0000",1598=> X"0000",1599=> X"0000",
                                        1600=> X"ffff",1601=> X"ffff",1602=> X"ff00",1603=> X"0000",1604=> X"0000",1605=> X"0000",1606=> X"0000",1607=> X"0000",1608=> X"8000",1609=> X"0000",1610=> X"0100",1611=> X"0000",1612=> X"0000",1613=> X"0000",1614=> X"0000",1615=> X"0000",1616=> X"8000",1617=> X"0000",1618=> X"0100",1619=> X"0000",1620=> X"0000",1621=> X"0000",1622=> X"0000",1623=> X"0000",1624=> X"8000",1625=> X"0000",1626=> X"0100",1627=> X"0000",1628=> X"0000",1629=> X"0000",1630=> X"0000",1631=> X"0000",1632=> X"8000",1633=> X"00f8",1634=> X"0100",1635=> X"0000",1636=> X"0000",1637=> X"0000",1638=> X"0000",1639=> X"0000",1640=> X"8000",1641=> X"018c",1642=> X"0100",1643=> X"0000",1644=> X"0000",1645=> X"0000",1646=> X"0000",1647=> X"0000",1648=> X"8000",1649=> X"0104",1650=> X"0100",1651=> X"0000",1652=> X"0000",1653=> X"0000",1654=> X"0000",1655=> X"0000",1656=> X"8000",1657=> X"0306",1658=> X"0100",1659=> X"0000",1660=> X"0000",1661=> X"0000",1662=> X"0000",1663=> X"0000",1664=> X"8000",1665=> X"0202",1666=> X"0100",1667=> X"0000",1668=> X"0000",1669=> X"0000",1670=> X"0000",1671=> X"0000",1672=> X"8000",1673=> X"1e02",1674=> X"0100",1675=> X"0000",1676=> X"0000",1677=> X"0000",1678=> X"0000",1679=> X"0000",1680=> X"8000",1681=> X"0202",1682=> X"0100",1683=> X"0000",1684=> X"0000",1685=> X"0000",1686=> X"0000",1687=> X"0000",1688=> X"8000",1689=> X"0202",1690=> X"0100",1691=> X"0000",1692=> X"0000",1693=> X"0000",1694=> X"0000",1695=> X"0000",1696=> X"8000",1697=> X"0202",1698=> X"0100",1699=> X"0000",1700=> X"0000",1701=> X"0000",1702=> X"0000",1703=> X"0000",1704=> X"8fff",1705=> X"e200",1706=> X"0100",1707=> X"0000",1708=> X"0000",1709=> X"0000",1710=> X"0000",1711=> X"0000",1712=> X"8000",1713=> X"2000",1714=> X"0100",1715=> X"0000",1716=> X"0000",1717=> X"0000",1718=> X"0000",1719=> X"0000",1720=> X"8000",1721=> X"2000",1722=> X"0700",1723=> X"0000",1724=> X"0000",1725=> X"0000",1726=> X"0000",1727=> X"0000",1728=> X"8000",1729=> X"2000",1730=> X"0100",1731=> X"0000",1732=> X"0000",1733=> X"0000",1734=> X"0000",1735=> X"0000",1736=> X"8000",1737=> X"2000",1738=> X"0100",1739=> X"0000",1740=> X"0000",1741=> X"0000",1742=> X"0000",1743=> X"0000",1744=> X"8000",1745=> X"2000",1746=> X"0100",1747=> X"0000",1748=> X"0000",1749=> X"0000",1750=> X"0000",1751=> X"0000",1752=> X"8000",1753=> X"2000",1754=> X"0100",1755=> X"0000",1756=> X"0000",1757=> X"0000",1758=> X"0000",1759=> X"0000",1760=> X"8000",1761=> X"2000",1762=> X"0100",1763=> X"0000",1764=> X"0000",1765=> X"0000",1766=> X"0000",1767=> X"0000",1768=> X"800f",1769=> X"fffc",1770=> X"0100",1771=> X"0000",1772=> X"0000",1773=> X"0000",1774=> X"0000",1775=> X"0000",1776=> X"8038",1777=> X"0000",1778=> X"0100",1779=> X"0000",1780=> X"0000",1781=> X"0000",1782=> X"0000",1783=> X"0000",1784=> X"8068",1785=> X"0000",1786=> X"0700",1787=> X"0000",1788=> X"0000",1789=> X"0000",1790=> X"0000",1791=> X"0000",1792=> X"80c8",1793=> X"0000",1794=> X"0100",1795=> X"0000",1796=> X"0000",1797=> X"0000",1798=> X"0000",1799=> X"0000",1800=> X"8188",1801=> X"0000",1802=> X"0100",1803=> X"0000",1804=> X"0000",1805=> X"0000",1806=> X"0000",1807=> X"0000",1808=> X"8308",1809=> X"0000",1810=> X"0100",1811=> X"0000",1812=> X"0000",1813=> X"0000",1814=> X"0000",1815=> X"0000",1816=> X"8608",1817=> X"0000",1818=> X"0100",1819=> X"0000",1820=> X"0000",1821=> X"0000",1822=> X"0000",1823=> X"0000",1824=> X"8c08",1825=> X"0000",1826=> X"0100",1827=> X"0000",1828=> X"0000",1829=> X"0000",1830=> X"0000",1831=> X"0000",1832=> X"ffff",1833=> X"ffff",1834=> X"ff00",1835=> X"0000",1836=> X"0000",1837=> X"0000",1838=> X"0000",1839=> X"0000",1840=> X"0000",1841=> X"0000",1842=> X"0000",1843=> X"0000",1844=> X"0000",1845=> X"0000",1846=> X"0000",1847=> X"0000",1848=> X"0000",1849=> X"0000",1850=> X"0000",1851=> X"0000",1852=> X"0000",1853=> X"0000",1854=> X"0000",1855=> X"0000",1856=> X"0000",1857=> X"0000",1858=> X"0000",1859=> X"0000",1860=> X"0000",1861=> X"0000",1862=> X"0000",1863=> X"0000",1864=> X"0000",1865=> X"0000",1866=> X"0000",1867=> X"0000",1868=> X"0000",1869=> X"0000",1870=> X"0000",1871=> X"0000",1872=> X"0000",1873=> X"0000",1874=> X"0000",1875=> X"0000",1876=> X"0000",1877=> X"0000",1878=> X"0000",1879=> X"0000",1880=> X"0000",1881=> X"0000",1882=> X"0000",1883=> X"0000",1884=> X"0000",1885=> X"0000",1886=> X"0000",1887=> X"0000",1888=> X"0000",1889=> X"0000",1890=> X"0000",1891=> X"0000",1892=> X"0000",1893=> X"0000",1894=> X"0000",1895=> X"0000",1896=> X"0000",1897=> X"0000",1898=> X"0000",1899=> X"0000",1900=> X"0000",1901=> X"0000",1902=> X"0000",1903=> X"0000",1904=> X"0000",1905=> X"0000",1906=> X"0000",1907=> X"0000",1908=> X"0000",1909=> X"0000",1910=> X"0000",1911=> X"0000",1912=> X"0000",1913=> X"0000",1914=> X"0000",1915=> X"0000",1916=> X"0000",1917=> X"0000",1918=> X"0000",1919=> X"0000",
                                      others=> X"0000");

    -- Micro memory
    type uMem_type is array (0 to 511) of STD_LOGIC_VECTOR(31 downto 0);
    constant uMem : uMem_type := (  0=>X"04100000",
                                    1=>X"03280000",
                                    2=>X"00000400",
                                    3=>X"0A540200",
                                    4=>X"04180000",
                                    5=>X"03500200",
                                    6=>X"04180000",
                                    7=>X"03100000",
                                    8=>X"03500200",
                                    9=>X"05A00600",
                                    10=>X"05100000",
                                    11=>X"0A300600",
                                    12=>X"15000000",
                                    13=>X"4A000000",
                                    14=>X"07A00600",
                                    15=>X"05400600",
                                    16=>X"00002A0F",
                                    17=>X"00000600",
                                    18=>X"0000220F",
                                    19=>X"00000600",
                                    20=>X"0000240F",
                                    21=>X"00000600",
                                    22=>X"00003816",
                                    23=>X"00000600",
                                    24=>X"1A000000",
                                    25=>X"55000600",
                                    26=>X"09100000",
                                    27=>X"04300000",
                                    28=>X"05420600",
                                    29=>X"00010000",
                                    30=>X"09100000",
                                    31=>X"03400600",
                                    32=>X"09100000",
                                    33=>X"0A320600",
                                    34=>X"00010000",
                                    35=>X"09100000",
                                    36=>X"03A00600",
                                    37=>X"05900600",
                                    38=>X"1A000000",
                                    39=>X"55000000",
                                    40=>X"07A00600",
                                    41=>X"05008000",
                                    42=>X"1A00342D",
                                    43=>X"D0004000",
                                    44=>X"0000322B",
                                    45=>X"07A00600",
                                    46=>X"05008000",
                                    47=>X"1A003432",
                                    48=>X"90004000",
                                    49=>X"00003230",
                                    50=>X"07A00600",
                                    51=>X"15000000",
                                    52=>X"6A000000",
                                    53=>X"07A00600",
                                    54=>X"15000000",
                                    55=>X"7A000000",
                                    56=>X"07A00600",
                                    57=>X"04180000",
                                    58=>X"13000000",
                                    59=>X"4A040000",
                                    60=>X"07100000",
                                    61=>X"03500200",
                                    62=>X"0000260F",
                                    63=>X"00000600",
                                    64=>X"0000280F",
                                    65=>X"00000600",
                                    66=>X"30000000",
                                    67=>X"55000000",
                                    68=>X"07A00600",
                                    69=>X"05008000",
                                    70=>X"00003846",
                                    71=>X"00007246",
                                    72=>X"00000600",
                                    511=>X"00003E00",
                                    others=> X"00000000");

    -- uPC
    signal uPC : STD_LOGIC_VECTOR(8 downto 0) := (others=>'0');
    signal SuPC : STD_LOGIC_VECTOR(8 downto 0) := (others=>'0');

    signal ctrlword : STD_LOGIC_VECTOR(31 downto 0) := X"00000000";
    alias cALU : STD_LOGIC_VECTOR(3 downto 0) is ctrlword(31 downto 28);
    alias cTB : STD_LOGIC_VECTOR(3 downto 0) is ctrlword(27 downto 24);
    alias cFB : STD_LOGIC_VECTOR(3 downto 0) is ctrlword(23 downto 20);
    alias cP : STD_LOGIC is ctrlword(19);
    alias cM : STD_LOGIC is ctrlword(18);
    alias cSP : STD_LOGIC_VECTOR(1 downto 0) is ctrlword(17 downto 16);
    alias cLC : STD_LOGIC_VECTOR(1 downto 0) is ctrlword(15 downto 14);
    alias cSEQ : STD_LOGIC_VECTOR(4 downto 0) is ctrlword(13 downto 9);
    alias cADR : STD_LOGIC_VECTOR(8 downto 0) is ctrlword(8 downto 0);

    type K1_type is array (0 to 63) of STD_LOGIC_VECTOR(8 downto 0);
    signal K1 : K1_type := (0=>"000001001", --MOVE
                            1=>"000001010", --STORE
                            2=>"000001100", --ADD
                            3=>"000001111", --BRA
                            4=>"000010000", --BCS
                            5=>"000010010", --BEQ
                            6=>"000010100", --BNE
                            7=>"000010110", --WVS
                            8=>"000011000", --CMP
                            9=>"000011010", --JSR
                            10=>"000011101", --RTS
                            11=>"000100000", --PUSH
                            12=>"000100010", --POP
                            13=>"000100101", --SSP
                            14=>"000100110", --SUB
                            15=>"000101001", --LSR
                            16=>"000101110", --LSL
                            17=>"000110011", --AND
                            18=>"000110110", --OR
                            19=>"000111110", --BMI
                            20=>"001000000", --BPL
                            21=>"001000010", --INV
                            22=>"001000101", --LWVS  
                            others=>"111111111"); --HULT

    type K2_type is array (0 to 3) of STD_LOGIC_VECTOR(8 downto 0);
    signal K2 : K2_type := (0=>"000000011", --reg-reg
                            1=>"000000100", --imm
                            2=>"000000110", --indir
                            3=>"000111001", --index
                            others=>"000000000");

    type gr_array is array (0 to 15) of STD_LOGIC_VECTOR(15 downto 0);
    signal rGR : gr_array := (others=> X"0000");

    signal tempGR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal tempPM : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal tempMM : STD_LOGIC_VECTOR(15 downto 0) := X"0000";


    ---------- DEBUG --------
    signal old_step : STD_LOGIC := '0';

begin
    ctrlword <= uMem(conv_integer(uPC));

    led_driver: leddriver port map (clk, rst, seg, an, led, rGR(2), rGR(5)(0) & rGR(4)(0) & "00000" & rGR(3)(0)); --rGR(2) 7-seg, rGR(3) leds
    --led_driver: leddriver port map (clk, rst, seg, an, led, rGR(2), rGR(5)(7 downto 0)); --rGR(2) 7-seg, rGR(3) leds
    alu_instance: alu port map(clk, cALU, rAR, databus, rAR, fC, fZ, fN, fO);
    

    -- *****************************
    -- * CONTROL UNIT              *
    -- *****************************
    process(clk) begin
        if rising_edge(clk) then
            
            -- rst
            if rst = '1' then
                rPC <= X"0000";
                uPC <= "000000000";
            else

                -- LC control
                case cLC is
                    when "01" => rLC <= rLC - 1;
                    when "10" => rLC <= databus(7 downto 0);
                    when "11" => rLC <= cADR(7 downto 0);
                    when others => null;
                end case;

                -- P control
                if cP = '1' then
                    rPC <= rPC + 1; 
                end if;

                -- SP control
                case cSP is
                    when "01" => rSP <= rSP + 1;
                    when "10" => rSP <= rSP - 1;
                    when others => null;
                end case;

                -- SEQ
                case cSEQ is
                    when "00000" => uPC <= uPC + 1;
                    when "00001" => uPC <= K1(conv_integer(rIR(15 downto 10)));
                    when "00010" => uPC <= K2(conv_integer(rIR(9 downto 8)));
                    when "00011" => uPC <= "000000000";
                    when "10000" => uPC <= cADR;
                    when "10001" => if fZ = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10010" => if fZ = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10011" => if fN = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10100" => if fN = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10101" => if fC = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10110" => if fC = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10111" => if fO = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11000" => if fO = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11001" => if fL = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11010" => if fL = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11011" => if fV = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11100" => if fV = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11101" => 
                        uPC <= cADR; 
                        SuPC <= uPC+1;
                    when "11110" => uPC <= SuPC;
                    when "11111" => null;
                    when others => null;
                end case;
                
                -- FROM BUS
                case cFB is
                    when "0001" => rASR <= databus;
                    when "0010" => rIR <= databus;
                    when "0011" => 
                        if (rASR(15) = '0') then
                            PrimMem(conv_integer(rASR)) <= databus;
                        elsif (rASR(15 downto 12) = X"9") then -- VR
                            vr_i <= databus;
                        end if;
                    when "0100" => rPC <= databus;
                    when "0101" => rDR <= databus;
                    when "0110" => null; -- can't write to uM
                    when "0111" => null; -- can't write to AR
                    when "1000" => rHR <= databus;
                    when "1001" => rSP <= databus;
                    when "1010" => 
                        if cM = '0' then 
                            rGR(conv_integer(rIR(7 downto 4))) <= databus;
                        else
                            rGR(conv_integer(rIR(3 downto 0))) <= databus;
                        end if;
                    when others => null;
                end case;
            end if;
        end if;
    end process;

    with rLC select
    fL <= '0' when X"00",
          '1' when others;

    --process(cFB, rASR, databus) begin
    process(clk) begin
        if rising_edge(clk) then
            if cFB = "0011" and rASR(15 downto 12) = X"9" then -- 9xxx address
                vr_we <= '1';
                --vr_i <= databus;
            else
                vr_we <= '0';
            end if;
        end if;
    end process;

    vr_addr <= rASR(4 downto 0);

    -- TO BUS
    with cTB select
    databus <= rASR when "0001",
                rIR when "0010",
                tempPM when "0011", -- PM/MM
                rPC when "0100",
                rDR when "0101",
                --uMem(conv_integer(uPC)) when "0110",
                rAR when "0111",
                rHR when "1000",
                rSP when "1001",
                tempGR when "1010",
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                --vr_o when "1011",
                X"0000" when others;

    -- PM/MemMap
    with rASR(15) select
    tempPM <= PrimMem(conv_integer(rASR)) when '0',
              tempMM when others;

    -- MemMap
    with rASR select
    tempMM <= "000000000000000" & up when X"8000",
              "000000000000000" & right when X"8001",
              "000000000000000" & down when X"8002",
              "000000000000000" & left when X"8003",
              X"00" & sw when X"8004",
              --X"00" & ledval when X"A000",
              --value when X"A001",
              vr_o when X"9000",vr_o when X"9001",vr_o when X"9002",vr_o when X"9003",
              vr_o when X"9004",vr_o when X"9005",vr_o when X"9006",vr_o when X"9007",
              vr_o when X"9008",vr_o when X"9009",vr_o when X"900A",vr_o when X"900B",
              vr_o when X"900C",vr_o when X"900D",vr_o when X"900E",vr_o when X"900F",
              vr_o when X"9010",vr_o when X"9011",vr_o when X"9012",vr_o when X"9013",
              vr_o when X"9014",vr_o when X"9015",vr_o when X"9016",vr_o when X"9017",
              vr_o when X"9018",vr_o when X"9019",vr_o when X"901A",vr_o when X"901B",
              vr_o when X"901C",vr_o when X"901D",vr_o when X"901E",vr_o when X"901F",
              X"EEEE" when others;

    -- M bit
    with cM select
    tempGR <= rGR(conv_integer(rIR(7 downto 4))) when '0',
              rGR(conv_integer(rIR(3 downto 0))) when others;

end cpu_one;
