library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity gpu is
    Port ( clk,rst : in  STD_LOGIC;
            vgaRed, vgaGreen: out STD_LOGIC_VECTOR (2 downto 0);
            vgaBlue : out STD_LOGIC_VECTOR (2 downto 1);
            Hsync,Vsync : out STD_LOGIC;
            vr_we : in STD_LOGIC;
            vr_addr: in STD_LOGIC_VECTOR(4 downto 0);
            vr_i: in STD_LOGIC_VECTOR(15 downto 0);
            vr_o: out STD_LOGIC_VECTOR(15 downto 0);
            fV: out STD_LOGIC);
end gpu;

architecture gpu_one of gpu is

    signal xctr,yctr : STD_LOGIC_VECTOR(11 downto 0) := "000000000000";
    alias xtile : STD_LOGIC_VECTOR(6 downto 0) is xctr(10 downto 4);
    alias ytile : STD_LOGIC_VECTOR(6 downto 0) is yctr(10 downto 4);
    alias tilexoff : STD_LOGIC_VECTOR(3 downto 0) is xctr(3 downto 0);
    alias tileyoff : STD_LOGIC_VECTOR(3 downto 0) is yctr(3 downto 0);
    signal hs : STD_LOGIC := '1';
    signal vs : STD_LOGIC := '1';
    signal pixel : STD_LOGIC_VECTOR(1 downto 0) := "00";
    signal video : STD_LOGIC_VECTOR(7 downto 0) := "00000000";
    alias red : STD_LOGIC_VECTOR(2 downto 0) is video(6 downto 4);
    alias green : STD_LOGIC_VECTOR(1 downto 0) is video(3 downto 2);
    alias blue : STD_LOGIC_VECTOR(1 downto 0) is video(1 downto 0);


    -- Tiles
    type pixel_data_type is array (0 to 255) of STD_LOGIC_VECTOR(7 downto 0);
    type tile_pixel_mem_type is array (0 to 31) of pixel_data_type;
    signal tile_pixel_mem : tile_pixel_mem_type := (
             0 => (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
             1 => (X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80"),
             2 => (X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80"),
             3 => (X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80"),
             4 => (X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"da",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
             5 => (X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90"),
             6 => (X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"da",X"da",X"da",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"ff",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"ff",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"ff",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"ff",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"c0",X"da",X"da",X"da",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"ff",X"c0",X"da",X"da",X"da",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"c0",X"da",X"da",X"da",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"ff",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"c0",X"da",X"da",X"da"),
             7 => (X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ea",X"da",X"ea",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ea",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da"),
             8 => (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"e0",X"e0",X"e0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"e0",X"e0",X"f0",X"e0",X"f0",X"e0",X"e0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"e0",X"f0",X"fd",X"fd",X"fd",X"f0",X"e0",X"f0",X"e0",X"00",X"00",X"00",X"00",X"00",X"00",X"e0",X"f0",X"fd",X"fd",X"f0",X"f0",X"f0",X"f0",X"e0",X"f0",X"e0",X"00",X"00",X"00",X"00",X"e0",X"f0",X"fd",X"fd",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"e0",X"00",X"00",X"00",X"e0",X"e0",X"fd",X"f0",X"f0",X"e0",X"f0",X"f0",X"e0",X"f0",X"e0",X"d0",X"e0",X"00",X"00",X"e0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"e0",X"f0",X"f0",X"f0",X"e0",X"f0",X"e0",X"00",X"e0",X"f0",X"f0",X"e0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"e0",X"d0",X"e0",X"e0",X"00",X"e0",X"f0",X"e0",X"f0",X"f0",X"e0",X"f0",X"f0",X"e0",X"f0",X"e0",X"f0",X"e0",X"d0",X"e0",X"00",X"00",X"e0",X"f0",X"e0",X"f0",X"f0",X"f0",X"f0",X"f0",X"e0",X"f0",X"e0",X"f0",X"e0",X"00",X"00",X"00",X"e0",X"e0",X"d0",X"e0",X"d0",X"e0",X"f0",X"e0",X"f0",X"e0",X"d0",X"e0",X"e0",X"00",X"00",X"00",X"00",X"e0",X"e0",X"f0",X"e0",X"f0",X"e0",X"d0",X"e0",X"f0",X"e0",X"e0",X"00",X"00",X"00",X"00",X"00",X"00",X"e0",X"e0",X"d0",X"e0",X"d0",X"e0",X"d0",X"e0",X"e0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"e0",X"e0",X"d0",X"e0",X"d0",X"e0",X"e0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"e0",X"e0",X"e0",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
             9 => (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"e8",X"e8",X"e8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"e8",X"e8",X"f8",X"f8",X"f8",X"e8",X"e8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"e8",X"f8",X"f8",X"fc",X"fc",X"fc",X"f8",X"f8",X"e8",X"00",X"00",X"00",X"00",X"00",X"00",X"e8",X"f8",X"f8",X"fc",X"fc",X"f8",X"f8",X"f8",X"f8",X"f8",X"e8",X"00",X"00",X"00",X"00",X"e8",X"f8",X"f8",X"fc",X"fc",X"f8",X"f8",X"e8",X"f8",X"f8",X"f8",X"f8",X"e8",X"00",X"00",X"00",X"e8",X"f8",X"fc",X"fc",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"e8",X"f8",X"e8",X"00",X"00",X"e8",X"f8",X"f8",X"fc",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"e8",X"00",X"e8",X"e8",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"e8",X"f8",X"f8",X"f8",X"f8",X"e8",X"e8",X"00",X"e8",X"f8",X"f8",X"f8",X"e8",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"e8",X"f8",X"e8",X"00",X"00",X"e8",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"f8",X"e8",X"f8",X"e8",X"00",X"00",X"00",X"e8",X"e8",X"f8",X"e8",X"f8",X"f8",X"f8",X"e8",X"f8",X"e8",X"f8",X"e8",X"e8",X"00",X"00",X"00",X"00",X"e8",X"e8",X"f8",X"e8",X"f8",X"e8",X"f8",X"e8",X"f8",X"e8",X"e8",X"00",X"00",X"00",X"00",X"00",X"00",X"e8",X"e8",X"f8",X"e8",X"f8",X"e8",X"f8",X"e8",X"e8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"e8",X"e8",X"f8",X"e8",X"f8",X"e8",X"e8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"e8",X"e8",X"e8",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
            10 => (X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"cf",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"df",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"ff",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"df",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80"),
            11 => (X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80"),
            12 => (X"da",X"da",X"c0",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"da",X"da",X"c0",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"da",X"da",X"c0",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"da",X"da",X"c0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"da",X"da",X"c0",X"80",X"ff",X"00",X"ff",X"00",X"ff",X"00",X"ff",X"00",X"ff",X"00",X"ff",X"00",X"da",X"da",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"da",X"da",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da"),
            13 => (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"ff",X"00",X"80",X"ff",X"00",X"ff",X"00",X"ff",X"00",X"ff",X"00",X"ff",X"00",X"ff",X"00",X"ff",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da"),
            14 => (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"ff",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"ff",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"ff",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"ff",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"ff",X"c0",X"da",X"da",X"da",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"c0",X"da",X"da",X"da",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"ff",X"c0",X"da",X"da",X"da",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"c0",X"da",X"da",X"da",X"80",X"ff",X"00",X"ff",X"00",X"ff",X"00",X"ff",X"00",X"ff",X"00",X"ff",X"c0",X"da",X"da",X"da",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"da",X"da",X"da",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"b0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da"),
            15 => (X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da"),
            16 => (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"8c",X"8c",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"9d",X"9d",X"9d",X"8c",X"9d",X"88",X"94",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"9d",X"9d",X"8c",X"a8",X"88",X"a8",X"88",X"89",X"88",X"00",X"00",X"00",X"00",X"00",X"88",X"9d",X"8c",X"88",X"a8",X"88",X"a8",X"94",X"a8",X"94",X"88",X"00",X"00",X"00",X"00",X"88",X"88",X"8c",X"a8",X"88",X"a8",X"94",X"a8",X"88",X"a8",X"94",X"88",X"89",X"00",X"00",X"00",X"88",X"88",X"89",X"88",X"a8",X"94",X"88",X"88",X"a8",X"89",X"88",X"94",X"88",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"a8",X"88",X"94",X"88",X"a8",X"94",X"94",X"94",X"00",X"00",X"00",X"00",X"89",X"88",X"88",X"89",X"88",X"a8",X"88",X"89",X"94",X"88",X"89",X"00",X"00",X"00",X"00",X"00",X"88",X"94",X"94",X"a8",X"a8",X"94",X"a8",X"88",X"94",X"89",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"89",X"94",X"a8",X"88",X"89",X"94",X"a8",X"94",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"a8",X"94",X"88",X"94",X"88",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"94",X"89",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
            17 => (X"00",X"00",X"00",X"00",X"00",X"00",X"8b",X"df",X"df",X"8b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"88",X"8b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"a8",X"88",X"8b",X"8b",X"8b",X"8b",X"88",X"8b",X"a8",X"a8",X"00",X"00",X"00",X"00",X"00",X"88",X"a8",X"a8",X"8b",X"8b",X"8b",X"b8",X"8b",X"a8",X"a8",X"88",X"a8",X"00",X"00",X"00",X"a8",X"a8",X"a8",X"8b",X"8b",X"8b",X"8b",X"88",X"a8",X"88",X"a8",X"a8",X"8b",X"a8",X"00",X"00",X"a8",X"88",X"8b",X"8b",X"8b",X"8b",X"8b",X"a8",X"88",X"a8",X"a8",X"8b",X"a8",X"a8",X"00",X"a8",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"a8",X"8b",X"8b",X"a8",X"8b",X"a8",X"a8",X"a8",X"e8",X"a8",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"c8",X"c8",X"8b",X"8b",X"a8",X"a8",X"e8",X"e8",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"c8",X"c8",X"c8",X"c8",X"c8",X"c8",X"e8",X"e8",X"e8",X"a8",X"a8",X"a8",X"8b",X"8b",X"8b",X"8b",X"b8",X"b8",X"b8",X"c8",X"c8",X"c8",X"c8",X"e8",X"e8",X"00",X"a8",X"88",X"8b",X"8b",X"8b",X"8b",X"8b",X"b8",X"b8",X"b8",X"8b",X"c8",X"c8",X"8b",X"00",X"00",X"a8",X"a8",X"8b",X"8b",X"8b",X"8b",X"8b",X"c8",X"b8",X"c8",X"8b",X"8b",X"8b",X"8b",X"00",X"00",X"00",X"a8",X"8b",X"8b",X"8b",X"8b",X"8b",X"c8",X"c8",X"c8",X"8b",X"8b",X"8b",X"00",X"00",X"00",X"00",X"00",X"a8",X"8b",X"8b",X"8b",X"8b",X"8b",X"c8",X"8b",X"8b",X"8b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"a8",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"8b",X"8b",X"8b",X"8b",X"00",X"00",X"00",X"00",X"00",X"00"),
            18 => (X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"ff",X"80",X"ff",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80"),
            19 => (X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"ff",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80"),
            20 => (X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da"),
            21 => (X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ea",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ea",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ea",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ea",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ea",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ea",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da"),
            22 => (X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ea",X"da",X"ea",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ea",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ea",X"da",X"ea",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da"),
            23 => (X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"c0",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"ff",X"da",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"c0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"c0",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"c0",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"a0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"ea",X"da",X"ea",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"ea",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"da",X"c0",X"c0",X"da",X"da",X"da",X"da",X"da",X"da",X"da"),
            24 => (X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"a4",X"a4",X"a4",X"a4",X"a4",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"a4",X"a0",X"a4",X"a4",X"a4",X"a0",X"a4",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"a4",X"a4",X"a4",X"a4",X"a4",X"a4",X"a4",X"80",X"80",X"80",X"00",X"00",X"80",X"94",X"94",X"80",X"80",X"a4",X"a4",X"a4",X"a4",X"a4",X"80",X"94",X"94",X"94",X"80",X"00",X"94",X"94",X"80",X"84",X"80",X"a4",X"80",X"a4",X"80",X"a4",X"80",X"80",X"94",X"94",X"94",X"80",X"94",X"80",X"84",X"84",X"80",X"a4",X"80",X"a4",X"80",X"a4",X"80",X"84",X"80",X"94",X"94",X"80",X"94",X"80",X"84",X"84",X"80",X"a4",X"80",X"a4",X"80",X"a4",X"80",X"84",X"80",X"94",X"94",X"80",X"94",X"80",X"84",X"84",X"84",X"80",X"84",X"80",X"84",X"80",X"84",X"84",X"80",X"94",X"94",X"80",X"94",X"80",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"80",X"94",X"94",X"80",X"94",X"94",X"80",X"84",X"84",X"84",X"00",X"00",X"84",X"84",X"84",X"80",X"94",X"94",X"80",X"00",X"94",X"94",X"94",X"80",X"84",X"00",X"00",X"00",X"00",X"84",X"80",X"94",X"94",X"94",X"80",X"00",X"80",X"94",X"00",X"00",X"80",X"80",X"00",X"00",X"80",X"80",X"00",X"00",X"94",X"80",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
            25 => (X"00",X"00",X"00",X"00",X"00",X"00",X"c2",X"d2",X"d2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"d2",X"d2",X"d2",X"d2",X"d2",X"d2",X"d2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"d2",X"c2",X"d2",X"f7",X"f7",X"f7",X"f7",X"d2",X"d2",X"00",X"00",X"00",X"00",X"00",X"00",X"d2",X"d2",X"f7",X"f7",X"f7",X"c2",X"d2",X"d2",X"d2",X"c2",X"d2",X"00",X"00",X"00",X"00",X"d2",X"f7",X"f7",X"f7",X"f7",X"d2",X"d2",X"d2",X"c2",X"d2",X"d2",X"d2",X"c2",X"00",X"00",X"00",X"d2",X"f7",X"f7",X"f7",X"d2",X"d2",X"d2",X"d2",X"d2",X"d2",X"c2",X"d2",X"c2",X"00",X"00",X"d2",X"d2",X"f7",X"c2",X"d2",X"d2",X"d2",X"c2",X"d2",X"d2",X"d2",X"d2",X"c2",X"d2",X"c2",X"00",X"c2",X"d2",X"d2",X"d2",X"d2",X"c2",X"d2",X"d2",X"d2",X"c2",X"d2",X"c2",X"d2",X"c2",X"c2",X"00",X"d2",X"d2",X"c2",X"d2",X"d2",X"d2",X"d2",X"d2",X"d2",X"d2",X"d2",X"d2",X"c2",X"d2",X"c2",X"00",X"00",X"c2",X"d2",X"c2",X"d2",X"c2",X"d2",X"d2",X"d2",X"c2",X"d2",X"c2",X"d2",X"c2",X"00",X"00",X"00",X"c2",X"c2",X"d2",X"c2",X"d2",X"c2",X"d2",X"c2",X"d2",X"c2",X"d2",X"c2",X"c2",X"00",X"00",X"00",X"00",X"c2",X"c2",X"d2",X"c2",X"d2",X"c2",X"d2",X"c2",X"d2",X"c2",X"c2",X"00",X"00",X"00",X"00",X"00",X"00",X"c2",X"c2",X"d2",X"c2",X"d2",X"c2",X"d2",X"c2",X"c2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"c2",X"c2",X"d2",X"c2",X"d2",X"c2",X"c2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"c2",X"c2",X"c2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
            26 => (X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"c0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"c0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"80",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"b0",X"c0",X"b0",X"c0",X"b0",X"c0",X"80",X"f0",X"b0",X"c0",X"b0",X"c0",X"b0",X"c0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"c0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"c0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"80",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"f5",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"f5",X"d0",X"f5",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"f5",X"d0",X"f5",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"b0",X"c0",X"b0",X"c0",X"b0",X"c0",X"80",X"f0",X"b0",X"c0",X"b0",X"c0",X"b0",X"c0",X"80"),
            27 => (X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"c0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"c0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"80",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"b0",X"c0",X"b0",X"c0",X"b0",X"c0",X"80",X"f0",X"b0",X"c0",X"b0",X"c0",X"b0",X"c0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"c0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"c0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"80",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"f5",X"d0",X"f5",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"f5",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"f5",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"b0",X"c0",X"b0",X"c0",X"b0",X"c0",X"80",X"f0",X"b0",X"c0",X"b0",X"c0",X"b0",X"c0",X"80"),
            28 => (X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"92",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"92",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"80",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"92",X"83",X"92",X"83",X"92",X"83",X"80",X"8b",X"92",X"83",X"92",X"83",X"92",X"83",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"92",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"92",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"80",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"92",X"83",X"92",X"83",X"92",X"83",X"80",X"8b",X"92",X"83",X"92",X"83",X"92",X"83",X"80"),
            29 => (X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"92",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"92",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"80",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"87",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"87",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"92",X"83",X"92",X"83",X"92",X"83",X"80",X"8b",X"92",X"87",X"92",X"87",X"92",X"87",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"92",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"92",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"80",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"8b",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"ea",X"87",X"ea",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"83",X"80",X"8b",X"87",X"87",X"ea",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"ea",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"83",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"87",X"87",X"87",X"87",X"87",X"92",X"80",X"8b",X"92",X"83",X"92",X"83",X"92",X"83",X"80",X"8b",X"92",X"83",X"92",X"83",X"92",X"83",X"80"),
            30 => (X"00",X"00",X"00",X"00",X"00",X"f0",X"f0",X"f0",X"f0",X"f0",X"00",X"00",X"fe",X"fe",X"fe",X"00",X"00",X"00",X"00",X"00",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"fe",X"fe",X"00",X"00",X"00",X"00",X"00",X"b4",X"b4",X"b4",X"fe",X"fe",X"80",X"fe",X"00",X"f0",X"f0",X"f0",X"00",X"00",X"00",X"00",X"b4",X"fe",X"b4",X"fe",X"fe",X"fe",X"80",X"fe",X"fe",X"fe",X"f0",X"f0",X"00",X"00",X"00",X"00",X"b4",X"fe",X"b4",X"b4",X"fe",X"fe",X"fe",X"80",X"fe",X"fe",X"fe",X"f0",X"00",X"00",X"00",X"00",X"b4",X"b4",X"fe",X"fe",X"fe",X"fe",X"80",X"80",X"80",X"80",X"f0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"fe",X"fe",X"fe",X"fe",X"fe",X"fe",X"fe",X"f0",X"f0",X"00",X"00",X"00",X"00",X"f0",X"f0",X"f0",X"f0",X"92",X"f0",X"f0",X"f0",X"92",X"f0",X"f0",X"00",X"00",X"b4",X"fe",X"fe",X"f0",X"f0",X"f0",X"f0",X"f0",X"82",X"f0",X"f0",X"f0",X"92",X"00",X"00",X"b4",X"b4",X"fe",X"fe",X"fe",X"f0",X"f0",X"f0",X"f0",X"82",X"82",X"82",X"82",X"fc",X"82",X"82",X"b4",X"b4",X"00",X"fe",X"00",X"00",X"92",X"f0",X"82",X"82",X"fc",X"82",X"82",X"82",X"82",X"82",X"b4",X"b4",X"00",X"00",X"b4",X"b4",X"b4",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"b4",X"b4",X"00",X"b4",X"b4",X"b4",X"82",X"82",X"82",X"82",X"82",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"b4",X"b4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
            31 => (X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"c0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"c0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"80",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"b0",X"c0",X"b0",X"c0",X"b0",X"c0",X"80",X"f0",X"b0",X"c0",X"b0",X"c0",X"b0",X"c0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"c0",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"c0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"80",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"c0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"d0",X"d0",X"d0",X"d0",X"d0",X"b0",X"80",X"f0",X"b0",X"c0",X"b0",X"c0",X"b0",X"c0",X"80",X"f0",X"b0",X"c0",X"b0",X"c0",X"b0",X"c0",X"80")

        --others => (others =>X"00") -- transparent
        );
    attribute ram_style: string;
    attribute ram_style of tile_pixel_mem : signal is "block";
    
    type sprite_pixel_mem_type is array(0 to 7) of pixel_data_type;
    constant sprite_pixel_mem : sprite_pixel_mem_type := (
        1 => (X"00",X"00",X"00",X"00",X"00",X"f0",X"f0",X"f0",X"f0",X"f0",X"00",X"00",X"fe",X"fe",X"fe",X"00",X"00",X"00",X"00",X"00",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"fe",X"fe",X"00",X"00",X"00",X"00",X"00",X"a0",X"a0",X"a0",X"fe",X"fe",X"80",X"fe",X"00",X"f0",X"f0",X"f0",X"00",X"00",X"00",X"00",X"a0",X"fe",X"a0",X"fe",X"fe",X"fe",X"80",X"fe",X"fe",X"fe",X"f0",X"f0",X"00",X"00",X"00",X"00",X"a0",X"fe",X"a0",X"a0",X"fe",X"fe",X"fe",X"80",X"fe",X"fe",X"fe",X"f0",X"00",X"00",X"00",X"00",X"a0",X"a0",X"fe",X"fe",X"fe",X"fe",X"80",X"80",X"80",X"80",X"f0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"fe",X"fe",X"fe",X"fe",X"fe",X"fe",X"fe",X"f0",X"f0",X"00",X"00",X"00",X"00",X"f0",X"f0",X"f0",X"f0",X"92",X"f0",X"f0",X"f0",X"92",X"f0",X"f0",X"00",X"00",X"a0",X"fe",X"fe",X"f0",X"f0",X"f0",X"f0",X"f0",X"92",X"f0",X"f0",X"f0",X"92",X"00",X"00",X"a0",X"a0",X"fe",X"fe",X"fe",X"f0",X"f0",X"f0",X"f0",X"92",X"92",X"92",X"92",X"ec",X"92",X"92",X"a0",X"a0",X"00",X"fe",X"00",X"00",X"92",X"f0",X"92",X"92",X"ec",X"92",X"92",X"92",X"92",X"92",X"a0",X"a0",X"00",X"00",X"a0",X"a0",X"a0",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"92",X"a0",X"a0",X"00",X"a0",X"a0",X"a0",X"92",X"92",X"92",X"92",X"92",X"92",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"a0",X"a0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),
        0 => (X"85",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"85",X"85",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"ec",X"83",X"85",X"85",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"83",X"83",X"85",X"85",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"83",X"83",X"85",X"85",X"80",X"80",X"ff",X"ff",X"ff",X"ff",X"ff",X"ff",X"ff",X"ff",X"80",X"80",X"83",X"83",X"85",X"85",X"80",X"80",X"ff",X"ff",X"ff",X"ff",X"ff",X"ff",X"ff",X"ff",X"80",X"80",X"83",X"83",X"85",X"85",X"80",X"80",X"ff",X"ff",X"80",X"80",X"80",X"80",X"ff",X"ff",X"80",X"80",X"83",X"83",X"85",X"85",X"80",X"80",X"ff",X"ff",X"80",X"80",X"80",X"80",X"ff",X"ff",X"80",X"80",X"83",X"83",X"85",X"85",X"80",X"80",X"ff",X"ff",X"80",X"80",X"80",X"80",X"ff",X"ff",X"80",X"80",X"83",X"83",X"85",X"85",X"80",X"80",X"ff",X"ff",X"80",X"80",X"80",X"80",X"ff",X"ff",X"80",X"80",X"83",X"83",X"85",X"85",X"80",X"80",X"ff",X"ff",X"ff",X"ff",X"ff",X"ff",X"ff",X"ff",X"80",X"80",X"83",X"83",X"85",X"85",X"80",X"80",X"ff",X"ff",X"ff",X"ff",X"ff",X"ff",X"ff",X"ff",X"80",X"80",X"83",X"83",X"85",X"85",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"83",X"83",X"85",X"85",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"83",X"83",X"85",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"83",X"83",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"f0",X"83"),
        others => (others =>X"F0")
    ); 

    type tile_mem_row_type is array(0 to 99) of STD_LOGIC_VECTOR(7 downto 0);
    type tile_mem_type is array(0 to 39) of tile_mem_row_type;

    constant layer0_mem : tile_mem_type := (
        0=> (X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 1=> (X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 2=> (X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 3=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 4=> (X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"1b",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 5=> (X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"04",X"05",X"06",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 6=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"16",X"0c",X"0d",X"0e",X"16",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 7=> (X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"15",X"15",X"16",X"15",X"16",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 8=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"04",X"05",X"05",X"05",X"05",X"05",X"06",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 9=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"1b",X"1a",X"1a",X"0c",X"0d",X"0d",X"0d",X"0d",X"0d",X"0e",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),10=> (X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"16",X"16",X"16",X"15",X"16",X"15",X"16",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),11=> (X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"04",X"05",X"05",X"05",X"05",X"05",X"06",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),12=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"0c",X"0d",X"0d",X"0d",X"0d",X"0d",X"0e",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),13=> (X"1a",X"00",X"00",X"00",X"1f",X"1f",X"1f",X"1a",X"1f",X"1f",X"1a",X"1a",X"1f",X"1f",X"1a",X"1a",X"1a",X"1b",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),14=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),15=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"1b",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),16=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),17=> (X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),18=> (X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),19=> (X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),20=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),21=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"1b",X"1f",X"1f",X"1b",X"1f",X"1a",X"1a",X"1f",X"1b",X"1b",X"1a",X"1b",X"1a",X"1a",X"1b",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),22=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"1a",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),23=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"1f",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"1b",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),24=> (X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"1b",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),25=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",X"1f",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),26=> (X"1a",X"00",X"00",X"00",X"00",X"00",X"1a",X"1a",X"00",X"00",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),27=> (X"1a",X"00",X"00",X"00",X"00",X"1a",X"1b",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),28=> (X"1b",X"00",X"00",X"00",X"1b",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"1b",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1a",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),29=> (X"1b",X"1b",X"1b",X"1a",X"1f",X"1f",X"1f",X"1a",X"1a",X"1f",X"1b",X"1b",X"1a",X"1f",X"1f",X"1b",X"1f",X"1f",X"1f",X"1a",X"1b",X"1f",X"1f",X"1b",X"1b",X"1b",X"1a",X"1b",X"1b",X"1b",X"1a",X"1f",X"1a",X"1a",X"1f",X"1a",X"1b",X"1a",X"1a",X"1f",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),30=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),31=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),32=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),33=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),34=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),35=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),36=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),37=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),38=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),39=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00")

);
    constant layer1_mem : tile_mem_type := (
        0=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 1=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 2=> (X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 3=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 4=> (X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"1d",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 5=> (X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"04",X"05",X"06",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 6=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"15",X"0c",X"0d",X"0e",X"16",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1e",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 7=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"16",X"16",X"15",X"15",X"15",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 8=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"04",X"05",X"05",X"05",X"05",X"05",X"06",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 9=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"0c",X"0d",X"0d",X"0d",X"0d",X"0d",X"0e",X"1d",X"1c",X"1c",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),10=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"16",X"16",X"15",X"16",X"15",X"16",X"16",X"1d",X"07",X"16",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),11=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"04",X"05",X"05",X"05",X"05",X"05",X"06",X"1c",X"07",X"15",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"1d",X"1d",X"0f",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),12=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"0c",X"0d",X"0d",X"0d",X"0d",X"0d",X"0e",X"1c",X"07",X"16",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"15",X"15",X"16",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),13=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"17",X"0f",X"17",X"1d",X"1c",X"1c",X"1d",X"1d",X"1c",X"1c",X"1c",X"1c",X"1c",X"1d",X"1d",X"1c",X"1c",X"04",X"05",X"06",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),14=> (X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"05",X"06",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"0c",X"0d",X"0e",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),15=> (X"1c",X"1c",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0c",X"0d",X"0e",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"0f",X"1c",X"1d",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),16=> (X"1c",X"00",X"1d",X"1c",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"15",X"14",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"04",X"05",X"06",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),17=> (X"1c",X"00",X"00",X"00",X"1d",X"1d",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"16",X"07",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"0c",X"0d",X"0e",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),18=> (X"1c",X"00",X"00",X"00",X"00",X"00",X"1c",X"1c",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"05",X"06",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"15",X"15",X"16",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),19=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"1c",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0c",X"0d",X"0e",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"1c",X"1c",X"0f",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),20=> (X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1c",X"1c",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"16",X"07",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"16",X"16",X"16",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),21=> (X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1d",X"1d",X"1d",X"1c",X"1c",X"1d",X"1c",X"1d",X"1d",X"1d",X"1d",X"1d",X"1d",X"1c",X"1d",X"1d",X"1c",X"1d",X"00",X"00",X"00",X"00",X"00",X"1d",X"04",X"05",X"06",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),22=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"06",X"1d",X"00",X"00",X"00",X"00",X"00",X"1c",X"0c",X"0d",X"0e",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),23=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0c",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0e",X"1c",X"00",X"00",X"00",X"00",X"00",X"1c",X"0f",X"1d",X"1d",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),24=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"16",X"16",X"15",X"16",X"16",X"16",X"15",X"15",X"16",X"15",X"16",X"15",X"15",X"15",X"15",X"1c",X"00",X"00",X"00",X"00",X"00",X"1c",X"04",X"05",X"06",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),25=> (X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"0f",X"1d",X"00",X"00",X"00",X"00",X"00",X"1d",X"0c",X"0d",X"0e",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),26=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"16",X"15",X"15",X"16",X"16",X"15",X"15",X"15",X"16",X"15",X"16",X"16",X"15",X"16",X"15",X"1c",X"00",X"00",X"00",X"00",X"00",X"1d",X"16",X"16",X"16",X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),27=> (X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"05",X"06",X"1c",X"00",X"00",X"00",X"00",X"00",X"1c",X"1d",X"1d",X"0f",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),28=> (X"1d",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0c",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0d",X"0e",X"1c",X"00",X"00",X"00",X"00",X"00",X"14",X"16",X"14",X"16",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),29=> (X"1c",X"1d",X"1c",X"1c",X"1d",X"1d",X"1c",X"1c",X"1c",X"1c",X"1d",X"1d",X"1c",X"1c",X"1c",X"1c",X"1c",X"1c",X"1c",X"1d",X"1d",X"1d",X"1d",X"1d",X"1d",X"1d",X"1d",X"1d",X"1c",X"1c",X"1d",X"1d",X"1d",X"1d",X"1c",X"1d",X"1c",X"1d",X"1c",X"1c",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),30=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),31=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),32=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),33=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),34=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),35=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),36=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),37=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),38=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),39=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00")
);
    
    constant layer2_mem : tile_mem_type := (
        0=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 1=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 2=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 3=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 4=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 5=> (X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00"), 6=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 7=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 8=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"), 9=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),10=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),11=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),12=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00"),13=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),14=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),15=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),16=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),17=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),18=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),19=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),20=> (X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00"),21=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),22=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),23=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),24=> (X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),25=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),26=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),27=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00"),28=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),29=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),30=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),31=> (X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),32=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),33=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),34=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),35=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),36=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00"),37=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),38=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"),39=> (X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00")
        --others => (others => X"00")
);

    constant layer3_mem : tile_mem_type := (
        0=> (X"13",X"01",X"03",X"0b",X"01",X"01",X"01",X"01",X"01",X"0b",X"01",X"13",X"01",X"01",X"02",X"01",X"12",X"13",X"0a",X"02",X"13",X"13",X"03",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"13",X"01",X"01",X"13",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"12",X"0b",X"0b",X"01",X"0a",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"13",X"01",X"13",X"01",X"03",X"01",X"01",X"13",X"01",X"13",X"01",X"13",X"01",X"0a",X"01",X"01",X"01",X"01",X"01",X"13",X"13",X"13",X"01",X"01",X"13",X"13",X"13",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"0b",X"12",X"0b",X"0b",X"02"), 1=> (X"01",X"01",X"01",X"02",X"12",X"0b",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"12",X"0a",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"03",X"13",X"01",X"01",X"13",X"01",X"03",X"01",X"01",X"01",X"01",X"12",X"02",X"01",X"01",X"01",X"02",X"13",X"01",X"02",X"01",X"01",X"03",X"01",X"0a",X"12",X"01",X"0a",X"01",X"0a",X"01",X"13",X"13",X"01",X"13",X"01",X"01",X"01",X"01",X"02",X"0a",X"01",X"01",X"01",X"13",X"13",X"01",X"01",X"02",X"01",X"02",X"0a",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"0a",X"0b",X"01",X"01",X"01",X"03",X"01",X"13",X"01"), 2=> (X"13",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"01",X"01",X"13",X"01",X"13",X"01",X"01",X"13",X"12",X"01",X"01",X"02",X"03",X"01",X"01",X"0b",X"13",X"02",X"0a",X"01",X"01",X"13",X"01",X"01",X"03",X"13",X"03",X"01",X"01",X"01",X"13",X"02",X"01",X"03",X"01",X"13",X"01",X"01",X"01",X"13",X"03",X"0b",X"0a",X"13",X"13",X"03",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"13",X"13",X"01",X"01",X"0a",X"13",X"02",X"01",X"02",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"02",X"01",X"13",X"01",X"0a",X"12",X"02",X"01",X"12",X"13",X"0b",X"01",X"0b",X"02"), 3=> (X"0b",X"01",X"01",X"01",X"13",X"13",X"01",X"0b",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"03",X"01",X"02",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"02",X"12",X"03",X"01",X"13",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"13",X"13",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"0b",X"01",X"01",X"01",X"01",X"01",X"03",X"02",X"02",X"01",X"13",X"01",X"12",X"01",X"13",X"01",X"01",X"01",X"13",X"0a",X"01",X"01",X"02",X"02",X"01",X"01",X"13",X"01",X"13",X"01",X"13",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"0b",X"01",X"12",X"01",X"01",X"02",X"01",X"01",X"01",X"02"), 4=> (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"03",X"01",X"0a",X"13",X"01",X"12",X"0a",X"01",X"01",X"01",X"0a",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"01",X"0b",X"01",X"01",X"01",X"0b",X"01",X"01",X"01",X"13",X"01",X"13",X"13",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"13",X"01",X"02",X"03",X"02",X"01",X"01",X"01",X"0a",X"02",X"01",X"03",X"12",X"01",X"02",X"0b"), 5=> (X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"02",X"13",X"03",X"0a",X"13",X"01",X"01",X"01",X"01",X"12",X"01",X"13",X"01",X"03",X"01",X"03",X"0a",X"13",X"0a",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"03",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"01",X"0a",X"0b",X"0b",X"01",X"03",X"03",X"12",X"01",X"0a",X"0b",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"01",X"02",X"02",X"01",X"01",X"03",X"13",X"01",X"13",X"13",X"01",X"13",X"13",X"01",X"01",X"01",X"01",X"12",X"01",X"13",X"01",X"01",X"01",X"13",X"01",X"02",X"12",X"0b",X"03"), 6=> (X"01",X"02",X"01",X"01",X"01",X"02",X"01",X"01",X"03",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"0a",X"02",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0b",X"03",X"01",X"12",X"13",X"01",X"12",X"0a",X"01",X"01",X"13",X"01",X"01",X"02",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"13",X"01",X"12",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"02",X"12",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"02",X"0a"), 7=> (X"0a",X"13",X"01",X"02",X"01",X"01",X"01",X"01",X"03",X"12",X"02",X"0b",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"0b",X"13",X"01",X"02",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"13",X"01",X"0a",X"13",X"0b",X"01",X"13",X"01",X"01",X"02",X"12",X"01",X"13",X"0a",X"12",X"01",X"12",X"0b",X"0b",X"01",X"02",X"13",X"13",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"13",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"13",X"01",X"01",X"01",X"01",X"01",X"13",X"13",X"01",X"13",X"01",X"13",X"01",X"02",X"01",X"01"), 8=> (X"01",X"0b",X"01",X"13",X"02",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"12",X"01",X"12",X"01",X"01",X"12",X"13",X"01",X"03",X"01",X"03",X"01",X"03",X"01",X"02",X"01",X"03",X"03",X"12",X"01",X"01",X"13",X"01",X"01",X"01",X"03",X"13",X"0b",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"02",X"12",X"13",X"02",X"01",X"01",X"0a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"13",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"13",X"13",X"01",X"01",X"01",X"01",X"12",X"01",X"13"), 9=> (X"12",X"01",X"02",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"0b",X"01",X"0b",X"02",X"03",X"0b",X"01",X"01",X"01",X"13",X"01",X"01",X"0b",X"0a",X"03",X"13",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"0b",X"01",X"13",X"03",X"01",X"01",X"13",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"0b",X"01",X"01",X"0a",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"13",X"13",X"01",X"0b",X"01",X"0b",X"01",X"02",X"01",X"01"),10=> (X"13",X"02",X"01",X"13",X"13",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"12",X"01",X"12",X"01",X"01",X"12",X"02",X"01",X"02",X"0a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"13",X"13",X"0a",X"03",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"03",X"01",X"01",X"01",X"0b",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"13",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"13",X"01"),11=> (X"13",X"01",X"13",X"13",X"01",X"01",X"01",X"01",X"13",X"01",X"13",X"01",X"01",X"01",X"02",X"0b",X"03",X"0a",X"01",X"01",X"12",X"03",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"12",X"03",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"13",X"01",X"01",X"01",X"0a",X"01",X"12",X"03",X"13",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"13"),12=> (X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"13",X"13",X"01",X"13",X"12",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"12",X"01",X"13",X"01",X"01",X"0b",X"12",X"0b",X"01",X"0b",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"13",X"01",X"13",X"13",X"01",X"13",X"13",X"01",X"13",X"13",X"13",X"01",X"0a",X"01",X"13",X"0a",X"01",X"01",X"01",X"02",X"01",X"13",X"0a",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0b",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01"),13=> (X"01",X"13",X"01",X"01",X"01",X"0b",X"03",X"02",X"0a",X"01",X"13",X"01",X"01",X"03",X"01",X"02",X"0b",X"01",X"12",X"01",X"0b",X"0a",X"02",X"01",X"01",X"01",X"02",X"0a",X"01",X"01",X"01",X"01",X"02",X"12",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"13",X"13",X"03",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"13",X"01",X"01",X"03",X"12",X"01",X"02",X"01",X"02",X"01",X"12",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"03",X"01",X"02",X"01",X"01",X"01",X"13",X"01",X"02",X"12",X"12",X"01",X"01",X"01",X"01"),14=> (X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"02",X"01",X"01",X"01",X"03",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"0b",X"01",X"13",X"13",X"01",X"0a",X"01",X"02",X"01",X"12",X"01",X"02",X"01",X"01",X"03",X"01",X"12",X"01",X"01",X"01",X"12",X"01",X"01",X"0b",X"01",X"01",X"01",X"01",X"03",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"0a",X"0a",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"02",X"12",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"12",X"02",X"01",X"01",X"01",X"13",X"01",X"01",X"02",X"0a",X"01",X"12",X"01",X"13",X"13",X"01",X"13"),15=> (X"01",X"01",X"12",X"0b",X"13",X"01",X"13",X"01",X"01",X"01",X"0a",X"01",X"01",X"13",X"01",X"0b",X"02",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"0a",X"01",X"13",X"01",X"01",X"01",X"01",X"0a",X"02",X"01",X"03",X"01",X"01",X"12",X"01",X"01",X"03",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"0a",X"01",X"13",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"03",X"12",X"01",X"01",X"0a",X"01",X"0a",X"0b",X"01",X"03",X"0a",X"02",X"01",X"13",X"01",X"13"),16=> (X"01",X"01",X"01",X"01",X"03",X"01",X"13",X"01",X"01",X"0b",X"01",X"0a",X"12",X"01",X"03",X"01",X"0b",X"03",X"01",X"01",X"01",X"0a",X"0a",X"12",X"01",X"02",X"0b",X"01",X"01",X"01",X"13",X"13",X"01",X"01",X"01",X"03",X"13",X"01",X"03",X"03",X"12",X"0a",X"03",X"01",X"01",X"01",X"0a",X"01",X"02",X"01",X"01",X"0b",X"01",X"13",X"0b",X"01",X"0a",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"0a",X"03",X"13",X"12",X"12",X"01",X"01",X"02",X"02",X"01",X"03",X"0b",X"01",X"01",X"0b",X"0a",X"13",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01"),17=> (X"01",X"03",X"01",X"01",X"0b",X"0b",X"01",X"03",X"13",X"01",X"12",X"13",X"0b",X"01",X"03",X"01",X"01",X"0a",X"0b",X"03",X"12",X"0b",X"01",X"01",X"01",X"0a",X"12",X"01",X"01",X"13",X"13",X"01",X"02",X"03",X"01",X"13",X"03",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"01",X"02",X"01",X"13",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"01",X"03",X"03",X"01",X"01",X"03",X"03",X"01",X"0b",X"01",X"0b",X"13",X"01",X"0a",X"01",X"0a",X"0a",X"13",X"01",X"13",X"01",X"01",X"01",X"13",X"01",X"0a",X"02",X"13",X"01",X"01",X"13",X"01"),18=> (X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"13",X"01",X"13",X"01",X"01",X"01",X"01",X"0a",X"02",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"02",X"01",X"02",X"01",X"02",X"13",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"02",X"03",X"13",X"01",X"01",X"12",X"01",X"02",X"02",X"01",X"01",X"0b",X"01",X"01",X"01",X"01",X"02",X"01",X"02",X"13",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"02",X"12",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"01"),19=> (X"12",X"13",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"13",X"01",X"13",X"01",X"13",X"13",X"01",X"13",X"0b",X"01",X"01",X"02",X"0a",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"12",X"13",X"13",X"01",X"13",X"01",X"01",X"01",X"13",X"13",X"01",X"13",X"01",X"01",X"01",X"13",X"01",X"13",X"13",X"01",X"13",X"13",X"01",X"01",X"02",X"03",X"01",X"01",X"01",X"01",X"02",X"01",X"03",X"02",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"03",X"01",X"01",X"01",X"13",X"01"),20=> (X"01",X"01",X"01",X"01",X"0b",X"03",X"01",X"01",X"01",X"13",X"01",X"13",X"01",X"01",X"01",X"01",X"02",X"01",X"0a",X"13",X"01",X"03",X"02",X"01",X"01",X"01",X"13",X"01",X"12",X"0a",X"01",X"0b",X"02",X"01",X"13",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"01",X"13",X"13",X"01",X"13",X"01",X"03",X"01",X"01",X"01",X"03",X"12",X"01",X"01",X"01",X"03",X"0a",X"01",X"01",X"01",X"01",X"0b",X"01",X"0a",X"01",X"01",X"13",X"0b",X"01",X"01",X"01",X"0a",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"03",X"01",X"01",X"01",X"13",X"0a",X"01",X"12"),21=> (X"01",X"0b",X"01",X"01",X"01",X"03",X"0a",X"01",X"01",X"01",X"01",X"01",X"13",X"13",X"01",X"01",X"0b",X"01",X"01",X"0a",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"13",X"01",X"0b",X"01",X"03",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"01",X"03",X"03",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"01",X"0a",X"01",X"0a",X"01",X"01",X"0b",X"01",X"03",X"01",X"01",X"01",X"03",X"0b",X"03",X"0b",X"0a",X"01",X"03",X"03",X"02",X"03",X"0a",X"03",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"02",X"01",X"01",X"02",X"03"),22=> (X"01",X"0b",X"01",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"0a",X"03",X"0b",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"13",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"01",X"13",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"03",X"12",X"03",X"13",X"02",X"13",X"01",X"01",X"13",X"01",X"13",X"01",X"01",X"13",X"02",X"02",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"13",X"01",X"02",X"12",X"01",X"01",X"13",X"13",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"02",X"01",X"02"),23=> (X"01",X"01",X"0b",X"01",X"01",X"0a",X"03",X"01",X"01",X"01",X"0b",X"01",X"02",X"01",X"01",X"01",X"03",X"02",X"01",X"01",X"03",X"01",X"01",X"01",X"0a",X"02",X"01",X"0a",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"03",X"01",X"01",X"01",X"01",X"01",X"0b",X"02",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"0b",X"02",X"01",X"01",X"13",X"13",X"13",X"13",X"01",X"01",X"13",X"02",X"0b",X"0a",X"0b",X"01",X"0b",X"0a",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"0a",X"01",X"01",X"01",X"13",X"01",X"03",X"02",X"01"),24=> (X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"12",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"12",X"12",X"13",X"0b",X"13",X"0b",X"01",X"01",X"01",X"01",X"0b",X"01",X"13",X"01",X"01",X"01",X"13",X"01",X"12",X"01",X"01",X"01",X"01",X"13",X"01",X"12",X"01",X"0a",X"13",X"0a",X"0b",X"01",X"01",X"01",X"01",X"03",X"01",X"13",X"01",X"01",X"01",X"01",X"0a",X"0b",X"01",X"01",X"0a",X"13",X"02",X"03",X"02",X"01",X"01",X"01",X"13",X"01",X"03",X"13",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"12",X"01",X"12",X"01",X"01",X"13",X"13",X"01",X"01",X"01"),25=> (X"01",X"03",X"02",X"02",X"0b",X"01",X"13",X"01",X"13",X"01",X"13",X"01",X"0b",X"01",X"01",X"03",X"01",X"13",X"12",X"0a",X"02",X"01",X"01",X"0b",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"0b",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"13",X"0a",X"01",X"01",X"02",X"01",X"01",X"01",X"0a",X"12",X"0a",X"13",X"01",X"13",X"01",X"01",X"01",X"13",X"13",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"12",X"01",X"03",X"01",X"01",X"02",X"12",X"01",X"01",X"03",X"0b",X"01",X"01",X"01",X"01",X"0b",X"01",X"01",X"01",X"0b",X"01",X"01",X"13",X"01",X"13",X"01",X"01",X"01"),26=> (X"01",X"01",X"12",X"12",X"0a",X"01",X"13",X"01",X"01",X"03",X"13",X"01",X"01",X"01",X"0b",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"02",X"12",X"01",X"01",X"12",X"13",X"02",X"01",X"01",X"12",X"0a",X"01",X"13",X"03",X"13",X"0b",X"01",X"13",X"01",X"02",X"02",X"01",X"03",X"13",X"01",X"01",X"01",X"0b",X"03",X"01",X"01",X"13",X"02",X"01",X"01",X"01",X"13",X"01",X"01",X"0b",X"01",X"01",X"02",X"01",X"0b",X"0a",X"01",X"01",X"01",X"01",X"13",X"13",X"01",X"01",X"13",X"12",X"13",X"01",X"0b",X"01",X"13",X"01",X"0b",X"0a",X"13"),27=> (X"01",X"0a",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"03",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"02",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"03",X"01",X"01",X"03",X"01",X"01",X"12",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"0a",X"12",X"03",X"03",X"0b",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"0a",X"0b",X"0b",X"02",X"01",X"02",X"13",X"02",X"01",X"13",X"13",X"01",X"02",X"03",X"03",X"01",X"01",X"01",X"01",X"12",X"0b",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"02",X"13",X"03",X"12",X"01",X"01",X"01"),28=> (X"01",X"13",X"12",X"01",X"01",X"0a",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"0b",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"0b",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"0b",X"01",X"01",X"01",X"03",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"13",X"12",X"0b",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"0a",X"01",X"01",X"03",X"03",X"13",X"02",X"01",X"0b",X"13",X"13",X"01",X"02",X"01",X"01",X"01",X"13",X"01",X"02",X"03",X"01",X"01",X"01",X"01",X"01",X"0a",X"0a",X"01",X"0b",X"01",X"0a",X"03",X"01",X"13",X"01",X"01",X"12",X"12",X"01",X"01",X"01",X"12"),29=> (X"12",X"03",X"01",X"03",X"01",X"0b",X"01",X"01",X"01",X"01",X"01",X"01",X"0b",X"02",X"12",X"0b",X"0a",X"02",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"03",X"02",X"01",X"01",X"02",X"12",X"0a",X"01",X"01",X"01",X"02",X"01",X"01",X"02",X"02",X"01",X"0a",X"01",X"01",X"01",X"03",X"01",X"02",X"01",X"01",X"01",X"03",X"12",X"13",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"01",X"13",X"03",X"01",X"13",X"01",X"01",X"12",X"01",X"01",X"01",X"01",X"13",X"01",X"13",X"01",X"01",X"01",X"01",X"0b",X"01",X"01",X"01",X"12",X"13",X"01",X"0a",X"13",X"01",X"01",X"12"),30=> (X"01",X"12",X"0a",X"01",X"01",X"01",X"0a",X"0b",X"0a",X"01",X"01",X"13",X"01",X"0a",X"01",X"0b",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"0a",X"01",X"01",X"0b",X"01",X"01",X"0a",X"01",X"13",X"01",X"01",X"03",X"0a",X"01",X"02",X"01",X"01",X"02",X"01",X"13",X"01",X"0b",X"01",X"01",X"01",X"13",X"01",X"01",X"03",X"01",X"02",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"13",X"01",X"13",X"01",X"01",X"13",X"01",X"0b",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"03",X"01",X"01",X"01",X"01",X"03",X"12",X"0b",X"12",X"13",X"02",X"03",X"01",X"01",X"13",X"01",X"01",X"03",X"03",X"03"),31=> (X"13",X"01",X"01",X"01",X"0b",X"02",X"0a",X"02",X"01",X"01",X"13",X"01",X"01",X"13",X"01",X"0b",X"13",X"01",X"01",X"01",X"01",X"0b",X"01",X"0b",X"13",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"02",X"01",X"01",X"01",X"13",X"01",X"01",X"02",X"12",X"01",X"01",X"13",X"13",X"01",X"01",X"0b",X"01",X"02",X"02",X"01",X"01",X"02",X"01",X"01",X"13",X"0a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"01",X"13",X"01",X"01",X"01",X"0a",X"01",X"12",X"13",X"0b",X"01",X"01",X"01",X"02",X"03",X"02",X"13"),32=> (X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"12",X"0a",X"01",X"01",X"13",X"01",X"02",X"02",X"0a",X"01",X"13",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"13",X"01",X"13",X"01",X"01",X"13",X"01",X"01",X"01",X"13",X"13",X"01",X"01",X"01",X"01",X"01",X"13",X"13",X"13",X"01",X"0b",X"13",X"13",X"01",X"01",X"01",X"0a",X"01",X"13",X"01",X"02",X"12",X"01",X"02",X"13",X"01",X"03",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"03",X"01",X"13",X"01"),33=> (X"12",X"01",X"01",X"03",X"12",X"01",X"01",X"01",X"13",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"0b",X"01",X"01",X"01",X"03",X"03",X"01",X"01",X"13",X"01",X"0b",X"02",X"13",X"01",X"13",X"01",X"01",X"01",X"01",X"03",X"01",X"13",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"13",X"01",X"13",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"12",X"01",X"12",X"01",X"0b",X"01",X"01",X"0a",X"02",X"01",X"0a",X"03",X"13",X"13",X"02",X"03",X"01",X"02",X"03",X"01",X"01",X"13",X"01",X"13",X"01",X"13",X"13",X"01",X"12",X"01",X"01",X"0a"),34=> (X"01",X"01",X"01",X"0b",X"03",X"01",X"13",X"01",X"01",X"01",X"13",X"13",X"13",X"01",X"0a",X"13",X"13",X"02",X"03",X"01",X"13",X"01",X"01",X"02",X"01",X"13",X"01",X"03",X"01",X"0a",X"01",X"01",X"01",X"01",X"01",X"13",X"03",X"13",X"0a",X"01",X"13",X"01",X"13",X"01",X"01",X"13",X"13",X"01",X"13",X"01",X"01",X"13",X"01",X"13",X"13",X"12",X"03",X"01",X"01",X"01",X"01",X"0b",X"03",X"01",X"01",X"01",X"01",X"0a",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"02",X"03",X"01",X"01",X"01",X"01",X"02",X"0b",X"0a",X"0a",X"0b",X"02",X"01",X"01",X"13",X"01",X"13",X"01",X"01",X"01",X"13",X"01",X"0b",X"02",X"12"),35=> (X"02",X"01",X"01",X"13",X"01",X"01",X"01",X"02",X"01",X"01",X"01",X"01",X"01",X"12",X"0b",X"01",X"01",X"01",X"01",X"02",X"01",X"0b",X"03",X"0b",X"02",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"01",X"13",X"01",X"03",X"03",X"01",X"01",X"0a",X"13",X"0a",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"13",X"01",X"0b",X"02",X"01",X"12",X"0b",X"01",X"01",X"01",X"12",X"02",X"01",X"01",X"0b",X"03",X"12",X"01",X"13",X"13",X"13",X"13",X"13",X"01",X"01",X"13",X"0b",X"01",X"01"),36=> (X"0a",X"01",X"01",X"01",X"0b",X"01",X"03",X"12",X"03",X"01",X"01",X"13",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"0a",X"03",X"12",X"03",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"01",X"13",X"0a",X"01",X"02",X"01",X"12",X"02",X"0a",X"01",X"01",X"01",X"01",X"01",X"03",X"02",X"02",X"13",X"03",X"0a",X"01",X"01",X"0a",X"03",X"01",X"01",X"0a",X"01",X"01",X"01",X"02",X"03",X"01",X"01",X"0a",X"01",X"01",X"01",X"01",X"0a",X"01",X"13",X"13",X"01",X"03",X"01",X"02",X"01",X"13",X"13",X"13",X"01",X"01",X"01",X"0b",X"01",X"13",X"01"),37=> (X"13",X"01",X"13",X"13",X"01",X"01",X"01",X"01",X"0a",X"13",X"01",X"01",X"13",X"01",X"01",X"01",X"01",X"02",X"03",X"13",X"13",X"01",X"13",X"01",X"13",X"0b",X"01",X"03",X"01",X"01",X"01",X"0b",X"01",X"0a",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0a",X"0a",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"13",X"13",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0b",X"01",X"13",X"01",X"01",X"01",X"01",X"01",X"13",X"12",X"01",X"01",X"02",X"01",X"01",X"13",X"01",X"03",X"01",X"0b",X"02",X"01",X"01",X"01",X"01",X"13",X"13",X"01",X"01",X"01",X"13",X"01"),38=> (X"03",X"01",X"13",X"01",X"0a",X"01",X"12",X"01",X"01",X"03",X"01",X"02",X"01",X"01",X"13",X"01",X"0a",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"02",X"0b",X"01",X"01",X"0a",X"01",X"01",X"03",X"01",X"01",X"13",X"01",X"0a",X"01",X"01",X"01",X"01",X"01",X"0b",X"03",X"01",X"01",X"01",X"01",X"12",X"03",X"01",X"0b",X"03",X"01",X"01",X"12",X"01",X"01",X"01",X"02",X"13",X"03",X"01",X"0b",X"13",X"13",X"01",X"01",X"01",X"13",X"01",X"13",X"13",X"01",X"01",X"01",X"0a",X"01",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"12",X"01",X"01",X"01",X"01",X"01",X"13",X"13",X"01",X"0b",X"01",X"01"),39=> (X"13",X"01",X"13",X"01",X"0b",X"03",X"03",X"01",X"13",X"01",X"03",X"02",X"13",X"01",X"0b",X"13",X"01",X"01",X"0b",X"0b",X"01",X"01",X"01",X"13",X"01",X"13",X"01",X"01",X"01",X"13",X"01",X"01",X"13",X"01",X"01",X"01",X"13",X"13",X"13",X"01",X"01",X"01",X"01",X"13",X"01",X"01",X"13",X"02",X"01",X"0b",X"03",X"13",X"01",X"13",X"01",X"01",X"13",X"01",X"02",X"03",X"01",X"01",X"01",X"0b",X"01",X"01",X"12",X"01",X"03",X"0a",X"01",X"13",X"01",X"13",X"13",X"01",X"01",X"13",X"01",X"02",X"0b",X"01",X"0a",X"01",X"01",X"13",X"01",X"01",X"02",X"13",X"01",X"01",X"13",X"13",X"13",X"13",X"01",X"01",X"01",X"01")
);

    signal current_tile0 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_tile1 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_tile2 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_tile3 : STD_LOGIC_VECTOR(7 downto 0) := X"00";


    signal current_pixel0 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_pixel1 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_pixel2 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_pixel3 : STD_LOGIC_VECTOR(7 downto 0) := X"00";


    signal current_sprite_pixel0 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_sprite_pixeL1 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_sprite_pixel2 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_sprite_pixel3 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_sprite_pixel4 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_sprite_pixel5 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_sprite_pixel6 : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal current_sprite_pixel7 : STD_LOGIC_VECTOR(7 downto 0) := X"00";

    type vr_array is array (0 to 31) of STD_LOGIC_VECTOR(15 downto 0);
    signal rVR : vr_array := (others=> X"0000"); --17=> X"0050", 18=> X"FFF0", 

    alias sprite0_x_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(0);
    alias sprite0_y_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(1);
    alias sprite1_x_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(2);
    alias sprite1_y_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(3);
    alias sprite2_x_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(4);
    alias sprite2_y_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(5);
    alias sprite3_x_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(6);
    alias sprite3_y_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(7);
    alias sprite4_x_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(8);
    alias sprite4_y_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(9);
    alias sprite5_x_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(10);
    alias sprite5_y_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(11);
    alias sprite6_x_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(12);
    alias sprite6_y_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(13);
    alias sprite7_x_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(14);
    alias sprite7_y_displacement : STD_LOGIC_VECTOR(15 downto 0) is rVR(15);

    alias x_displacement0 : STD_LOGIC_VECTOR(15 downto 0) is rVR(16);
    alias y_displacement0 : STD_LOGIC_VECTOR(15 downto 0) is rVR(17);
    alias x_displacement1 : STD_LOGIC_VECTOR(15 downto 0) is rVR(18);
    alias y_displacement1 : STD_LOGIC_VECTOR(15 downto 0) is rVR(19);
    alias x_displacement2 : STD_LOGIC_VECTOR(15 downto 0) is rVR(20);
    alias y_displacement2 : STD_LOGIC_VECTOR(15 downto 0) is rVR(21);
    alias x_displacement3 : STD_LOGIC_VECTOR(15 downto 0) is rVR(22);
    alias y_displacement3 : STD_LOGIC_VECTOR(15 downto 0) is rVR(23);

    alias sprite_0_layer : STD_LOGIC_VECTOR(1 downto 0) is rVR(26)(15 downto 14);
    alias sprite_1_layer : STD_LOGIC_VECTOR(1 downto 0) is rVR(26)(13 downto 12);
    alias sprite_2_layer : STD_LOGIC_VECTOR(1 downto 0) is rVR(26)(11 downto 10);
    alias sprite_3_layer : STD_LOGIC_VECTOR(1 downto 0) is rVR(26)(9 downto 8);
    alias sprite_4_layer : STD_LOGIC_VECTOR(1 downto 0) is rVR(26)(7 downto 6);
    alias sprite_5_layer : STD_LOGIC_VECTOR(1 downto 0) is rVR(26)(5 downto 4);
    alias sprite_6_layer : STD_LOGIC_VECTOR(1 downto 0) is rVR(26)(3 downto 2);
    alias sprite_7_layer : STD_LOGIC_VECTOR(1 downto 0) is rVR(26)(1 downto 0);

    signal counter : STD_LOGIC_VECTOR(23 downto 0) := "000000000000000000000000";

    signal tilepix_addra : STD_LOGIC_VECTOR(4 downto 0) := "00000";
    signal tilepix_addrb : STD_LOGIC_VECTOR(4 downto 0) := "00000";
    signal tilepix_subaddra : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal tilepix_subaddrb : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal tilepix_dataina : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal tilepix_datainb : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal tilepix_datauta : STD_LOGIC_VECTOR(7 downto 0) := X"00";
    signal tilepix_datautb : STD_LOGIC_VECTOR(7 downto 0) := X"00";
begin
    
    --process(vr_i, vr_we, vr_addr, rst, rVR) begin
    process(clk) begin
        if rising_edge(clk) then
            if rst='1' then
                rVR <= (others=> X"0000");
            else
                if vr_we = '1' then
                    rVR(conv_integer(vr_addr)) <= vr_i;
                end if;
                vr_o <= rVR(conv_integer(vr_addr));
            end if;
        end if;
    end process;


    -- Tile pixel access
    process(clk) begin
        if rising_edge(clk) then
            tilepix_datauta <= tile_pixel_mem(conv_integer(tilepix_addra))(conv_integer(tilepix_subaddra));
            tilepix_datautb <= tile_pixel_mem(conv_integer(tilepix_addrb))(conv_integer(tilepix_subaddrb));
        end if;
    end process;

    -- Pixel clock
    process(clk) begin
     if rising_edge(clk) then
       if rst='1' then
         pixel <= "00";
       else
         pixel <= pixel + 1;
       end if;
     end if;
  end process;

  process(clk) begin
    if rising_edge(clk) then
      if rst='1' then
         xctr <= "000000000000";
      elsif pixel=3 then
       if xctr=799 then
         xctr <= "000000000000";
       else
         xctr <= xctr + 1;
       end if;
      end if;

      if xctr=656 then -- 688
        hs <= '0';
      elsif xctr=752 then -- 784
        hs <= '1';
      end if;
    end if;
  end process;

  process(clk) begin
    if rising_edge(clk) then
      if rst='1' then
        yctr <= "000000000000";
      elsif xctr=799 and pixel=0 then
       if yctr=520 then
         yctr <= "000000000000";
       else
         yctr <= yctr + 1;
       end if;

       if yctr=490 then -- 509
         vs <= '0';
       elsif  yctr=492 then --511
         vs <= '1';
       end if;
      end if;
    end if;
  end process;
  Hsync <= hs;
  Vsync <= vs;

  process(clk) begin
    if rising_edge(clk) then
        if yctr = 480 and xctr = 0 and pixel = "00" then
            fV <= '1';
        else
            fV <= '0'; -- Should be 0, debug
        end if;
    end if;
  end process;
     

  process(clk) begin
    if rising_edge(clk) then
        if yctr<479 and xctr<639 then
            if pixel = "00" then

                --
                -- Start of checking the current tiles
                --
                if xctr - x_displacement0 > 1599 or yctr - y_displacement0 > 639 then
                    current_tile0 <= X"00";
                elsif x_displacement0(3 downto 0) <= tilexoff and y_displacement0(3 downto 0) <= tileyoff  then 
                    current_tile0 <= layer0_mem(conv_integer(ytile) - conv_integer(y_displacement0(10 downto 4)))
                                               (conv_integer(xtile) - conv_integer(x_displacement0(10 downto 4)));
                elsif x_displacement0(3 downto 0) <= tilexoff then
                    current_tile0 <= layer0_mem(conv_integer(ytile) - conv_integer(y_displacement0(10 downto 4) + 1))
                                               (conv_integer(xtile) - conv_integer(x_displacement0(10 downto 4)));
                elsif y_displacement0(3 downto 0) <= tileyoff then
                    current_tile0 <= layer0_mem(conv_integer(ytile) - conv_integer(y_displacement0(10 downto 4)))
                                               (conv_integer(xtile) - conv_integer(x_displacement0(10 downto 4) + 1));
                else
                    current_tile0 <= layer0_mem(conv_integer(ytile) - conv_integer(y_displacement0(10 downto 4) + 1))
                                               (conv_integer(xtile) - conv_integer(x_displacement0(10 downto 4) + 1));
                end if;
                if xctr - x_displacement1 > 1599 or yctr - y_displacement1 > 639 then
                    current_tile1 <= X"00";
                elsif x_displacement1(3 downto 0) <= tilexoff and y_displacement1(3 downto 0) <= tileyoff  then 
                    current_tile1 <= layer1_mem(conv_integer(ytile) - conv_integer(y_displacement1(10 downto 4)))
                                               (conv_integer(xtile) - conv_integer(x_displacement1(10 downto 4)));
                elsif x_displacement1(3 downto 0) <= tilexoff then
                    current_tile1 <= layer1_mem(conv_integer(ytile) - conv_integer(y_displacement1(10 downto 4) + 1))
                                               (conv_integer(xtile) - conv_integer(x_displacement1(10 downto 4)));
                elsif y_displacement1(3 downto 0) <= tileyoff then
                    current_tile1 <= layer1_mem(conv_integer(ytile) - conv_integer(y_displacement1(10 downto 4)))
                                               (conv_integer(xtile) - conv_integer(x_displacement1(10 downto 4) + 1));
                else
                    current_tile1 <= layer1_mem(conv_integer(ytile) - conv_integer(y_displacement1(10 downto 4) + 1))
                                               (conv_integer(xtile) - conv_integer(x_displacement1(10 downto 4) + 1));
                end if;


                
            elsif pixel = "01" then --tile_pixel 0 and 1

                if xctr - x_displacement2 > 1599 or yctr - y_displacement2 > 639 then
                    current_tile2 <= X"00";
                elsif x_displacement2(3 downto 0) <= tilexoff and y_displacement2(3 downto 0) <= tileyoff  then 
                    current_tile2 <= layer2_mem(conv_integer(ytile) - conv_integer(y_displacement2(10 downto 4)))
                                               (conv_integer(xtile) - conv_integer(x_displacement2(10 downto 4)));
                elsif x_displacement2(3 downto 0) <= tilexoff then
                    current_tile2 <= layer2_mem(conv_integer(ytile) - conv_integer(y_displacement2(10 downto 4) + 1))
                                               (conv_integer(xtile) - conv_integer(x_displacement2(10 downto 4)));
                elsif y_displacement2(3 downto 0) <= tileyoff then
                    current_tile2 <= layer2_mem(conv_integer(ytile) - conv_integer(y_displacement2(10 downto 4)))
                                               (conv_integer(xtile) - conv_integer(x_displacement2(10 downto 4) + 1));
                else
                    current_tile2 <= layer2_mem(conv_integer(ytile) - conv_integer(y_displacement2(10 downto 4) + 1))
                                               (conv_integer(xtile) - conv_integer(x_displacement2(10 downto 4) + 1));
                end if;
                if xctr - x_displacement3 > 1599 or yctr - y_displacement3 > 639 then
                    current_tile3 <= X"00";
                elsif x_displacement3(3 downto 0) <= tilexoff and y_displacement3(3 downto 0) <= tileyoff  then 
                    current_tile3 <= layer3_mem(conv_integer(ytile) - conv_integer(y_displacement3(10 downto 4)))
                                               (conv_integer(xtile) - conv_integer(x_displacement3(10 downto 4)));
                elsif x_displacement3(3 downto 0) <= tilexoff then
                    current_tile3 <= layer3_mem(conv_integer(ytile) - conv_integer(y_displacement3(10 downto 4) + 1))
                                               (conv_integer(xtile) - conv_integer(x_displacement3(10 downto 4)));
                elsif y_displacement3(3 downto 0) <= tileyoff then
                    current_tile3 <= layer3_mem(conv_integer(ytile) - conv_integer(y_displacement3(10 downto 4)))
                                               (conv_integer(xtile) - conv_integer(x_displacement3(10 downto 4) + 1));
                else
                    current_tile3 <= layer3_mem(conv_integer(ytile) - conv_integer(y_displacement3(10 downto 4) + 1))
                                               (conv_integer(xtile) - conv_integer(x_displacement3(10 downto 4) + 1));
                end if;


                current_pixel0 <= tile_pixel_mem(conv_integer(current_tile0(4 downto 0)))(conv_integer((tileyoff - y_displacement0(3 downto 0)) & 
                                                                                                       (tilexoff - x_displacement0(3 downto 0))));
                current_pixel1 <= tile_pixel_mem(conv_integer(current_tile1(4 downto 0)))(conv_integer((tileyoff - y_displacement1(3 downto 0)) &
                                                                                                       (tilexoff - x_displacement1(3 downto 0))));
            elsif pixel = "10" then --sprite pixels and tile_pixel 2 and 3

                current_pixel2 <= tile_pixel_mem(conv_integer(current_tile2(4 downto 0)))(conv_integer((tileyoff - y_displacement2(3 downto 0)) &
                                                                                                       (tilexoff - x_displacement2(3 downto 0))));
                current_pixel3 <= tile_pixel_mem(conv_integer(current_tile3(4 downto 0)))(conv_integer((tileyoff - y_displacement3(3 downto 0)) &
                                                                                                       (tilexoff - x_displacement3(3 downto 0))));

                --
                -- Check sprite pixels
                --
                if xctr(11 downto 0) >= sprite0_x_displacement(15 downto 0) and xctr(11 downto 0) < sprite0_x_displacement(15 downto 0) + 16 and 
                   yctr(11 downto 0) >= sprite0_y_displacement(15 downto 0) and yctr(11 downto 0) < sprite0_y_displacement(15 downto 0) + 16 then
                    current_sprite_pixel0 <= sprite_pixel_mem(conv_integer(rVR(24)(15 downto 12)))(conv_integer((tileyoff - sprite0_y_displacement(3 downto 0)) & 
                                                                                                                (tilexoff - sprite0_x_displacement(3 downto 0))));
                else current_sprite_pixel0 <= X"00"; end if;
                if xctr(11 downto 0) >= sprite1_x_displacement(15 downto 0) and xctr(11 downto 0) < sprite1_x_displacement(15 downto 0) + 16 and 
                   yctr(11 downto 0) >= sprite1_y_displacement(15 downto 0) and yctr(11 downto 0) < sprite1_y_displacement(15 downto 0) + 16 then
                    current_sprite_pixel1 <= sprite_pixel_mem(conv_integer(rVR(24)(11 downto 8)))(conv_integer((tileyoff - sprite1_y_displacement(3 downto 0)) & 
                                                                                                               (tilexoff - sprite1_x_displacement(3 downto 0))));
                else current_sprite_pixel1 <= X"00"; end if;
                if xctr(11 downto 0) >= sprite2_x_displacement(15 downto 0) and xctr(11 downto 0) < sprite2_x_displacement(15 downto 0) + 16 and 
                   yctr(11 downto 0) >= sprite2_y_displacement(15 downto 0) and yctr(11 downto 0) < sprite2_y_displacement(15 downto 0) + 16 then
                    current_sprite_pixel2 <= sprite_pixel_mem(conv_integer(rVR(24)(7 downto 4)))(conv_integer((tileyoff - sprite2_y_displacement(3 downto 0)) & 
                                                                                                              (tilexoff - sprite2_x_displacement(3 downto 0))));
                else current_sprite_pixel2 <= X"00"; end if;
                if xctr(11 downto 0) >= sprite3_x_displacement(15 downto 0) and xctr(11 downto 0) < sprite3_x_displacement(15 downto 0) + 16 and 
                   yctr(11 downto 0) >= sprite3_y_displacement(15 downto 0) and yctr(11 downto 0) < sprite3_y_displacement(15 downto 0) + 16 then
                    current_sprite_pixel3 <= sprite_pixel_mem(conv_integer(rVR(24)(3 downto 0)))(conv_integer((tileyoff - sprite3_y_displacement(3 downto 0)) & 
                                                                                                              (tilexoff - sprite3_x_displacement(3 downto 0))));
                else current_sprite_pixel3 <= X"00"; end if;
                if xctr(11 downto 0) >= sprite4_x_displacement(15 downto 0) and xctr(11 downto 0) < sprite4_x_displacement(15 downto 0) + 16 and 
                   yctr(11 downto 0) >= sprite4_y_displacement(15 downto 0) and yctr(11 downto 0) < sprite4_y_displacement(15 downto 0) + 16 then
                    current_sprite_pixel4 <= sprite_pixel_mem(conv_integer(rVR(25)(15 downto 12)))(conv_integer((tileyoff - sprite4_y_displacement(3 downto 0)) & 
                                                                                                                (tilexoff - sprite4_x_displacement(3 downto 0))));
                else current_sprite_pixel4 <= X"00"; end if;
                if xctr(11 downto 0) >= sprite5_x_displacement(15 downto 0) and xctr(11 downto 0) < sprite5_x_displacement(15 downto 0) + 16 and 
                   yctr(11 downto 0) >= sprite5_y_displacement(15 downto 0) and yctr(11 downto 0) < sprite5_y_displacement(15 downto 0) + 16 then
                    current_sprite_pixel5 <= sprite_pixel_mem(conv_integer(rVR(25)(11 downto 8)))(conv_integer((tileyoff - sprite5_y_displacement(3 downto 0)) & 
                                                                                                               (tilexoff - sprite5_x_displacement(3 downto 0))));
                else current_sprite_pixel5 <= X"00"; end if;
                if xctr(11 downto 0) >= sprite6_x_displacement(15 downto 0) and xctr(11 downto 0) < sprite6_x_displacement(15 downto 0) + 16 and 
                   yctr(11 downto 0) >= sprite6_y_displacement(15 downto 0) and yctr(11 downto 0) < sprite6_y_displacement(15 downto 0) + 16 then
                    current_sprite_pixel6 <= sprite_pixel_mem(conv_integer(rVR(25)(11 downto 4)))(conv_integer((tileyoff - sprite6_y_displacement(3 downto 0)) & 
                                                                                                               (tilexoff - sprite6_x_displacement(3 downto 0))));
                else current_sprite_pixel6 <= X"00"; end if;
                if xctr(11 downto 0) >= sprite7_x_displacement(15 downto 0) and xctr(11 downto 0) < sprite7_x_displacement(15 downto 0) + 16 and 
                   yctr(11 downto 0) >= sprite7_y_displacement(15 downto 0) and yctr(11 downto 0) < sprite7_y_displacement(15 downto 0) + 16 then
                    current_sprite_pixel7 <= sprite_pixel_mem(conv_integer(rVR(25)(3 downto 0)))(conv_integer((tileyoff - sprite7_y_displacement(3 downto 0)) & 
                                                                                                              (tilexoff - sprite7_x_displacement(3 downto 0))));
                else current_sprite_pixel7 <= X"00"; end if;

            elsif pixel = "11" then --val av pixel
                if    sprite_0_layer = "00" and current_sprite_pixel0(7) = '1' then video <= current_sprite_pixel0; 
                elsif sprite_1_layer = "00" and current_sprite_pixel1(7) = '1' then video <= current_sprite_pixel1; 
                elsif sprite_2_layer = "00" and current_sprite_pixel2(7) = '1' then video <= current_sprite_pixel2; 
                elsif sprite_3_layer = "00" and current_sprite_pixel3(7) = '1' then video <= current_sprite_pixel3; 
                elsif sprite_4_layer = "00" and current_sprite_pixel4(7) = '1' then video <= current_sprite_pixel4; 
                elsif sprite_5_layer = "00" and current_sprite_pixel5(7) = '1' then video <= current_sprite_pixel5; 
                elsif sprite_6_layer = "00" and current_sprite_pixel6(7) = '1' then video <= current_sprite_pixel6; 
                elsif sprite_7_layer = "00" and current_sprite_pixel7(7) = '1' then video <= current_sprite_pixel7; 
                elsif current_pixel0(7) = '1' then video <= current_pixel0;
                elsif sprite_0_layer = "01" and current_sprite_pixel0(7) = '1' then video <= current_sprite_pixel0; 
                elsif sprite_1_layer = "01" and current_sprite_pixel1(7) = '1' then video <= current_sprite_pixel1; 
                elsif sprite_2_layer = "01" and current_sprite_pixel2(7) = '1' then video <= current_sprite_pixel2; 
                elsif sprite_3_layer = "01" and current_sprite_pixel3(7) = '1' then video <= current_sprite_pixel3; 
                elsif sprite_4_layer = "01" and current_sprite_pixel4(7) = '1' then video <= current_sprite_pixel4; 
                elsif sprite_5_layer = "01" and current_sprite_pixel5(7) = '1' then video <= current_sprite_pixel5; 
                elsif sprite_6_layer = "01" and current_sprite_pixel6(7) = '1' then video <= current_sprite_pixel6; 
                elsif sprite_7_layer = "01" and current_sprite_pixel7(7) = '1' then video <= current_sprite_pixel7; 
                elsif current_pixel1(7) = '1' then video <= current_pixel1;
                elsif sprite_0_layer = "10" and current_sprite_pixel0(7) = '1' then video <= current_sprite_pixel0; 
                elsif sprite_1_layer = "10" and current_sprite_pixel1(7) = '1' then video <= current_sprite_pixel1; 
                elsif sprite_2_layer = "10" and current_sprite_pixel2(7) = '1' then video <= current_sprite_pixel2; 
                elsif sprite_3_layer = "10" and current_sprite_pixel3(7) = '1' then video <= current_sprite_pixel3; 
                elsif sprite_4_layer = "10" and current_sprite_pixel4(7) = '1' then video <= current_sprite_pixel4; 
                elsif sprite_5_layer = "10" and current_sprite_pixel5(7) = '1' then video <= current_sprite_pixel5; 
                elsif sprite_6_layer = "10" and current_sprite_pixel6(7) = '1' then video <= current_sprite_pixel6; 
                elsif sprite_7_layer = "10" and current_sprite_pixel7(7) = '1' then video <= current_sprite_pixel7; 
                elsif current_pixel2(7) = '1' then video <= current_pixel2;
                elsif sprite_0_layer = "11" and current_sprite_pixel0(7) = '1' then video <= current_sprite_pixel0; 
                elsif sprite_1_layer = "11" and current_sprite_pixel1(7) = '1' then video <= current_sprite_pixel1; 
                elsif sprite_2_layer = "11" and current_sprite_pixel2(7) = '1' then video <= current_sprite_pixel2; 
                elsif sprite_3_layer = "11" and current_sprite_pixel3(7) = '1' then video <= current_sprite_pixel3; 
                elsif sprite_4_layer = "11" and current_sprite_pixel4(7) = '1' then video <= current_sprite_pixel4; 
                elsif sprite_5_layer = "11" and current_sprite_pixel5(7) = '1' then video <= current_sprite_pixel5; 
                elsif sprite_6_layer = "11" and current_sprite_pixel6(7) = '1' then video <= current_sprite_pixel6; 
                elsif sprite_7_layer = "11" and current_sprite_pixel7(7) = '1' then video <= current_sprite_pixel7; 
                else video <= current_pixel3;
                end if;
            end if;
        else
          video <= "00000000";
        end if;
    end if;
  end process;

  vgaRed(2 downto 0) <= (red);
  vgaGreen(2 downto 0) <= (green & '0');
  vgaBlue(2 downto 1) <= (blue);


end gpu_one;
