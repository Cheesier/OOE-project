library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity alu is
    Port (  clk : in STD_LOGIC;
            op : in STD_LOGIC_VECTOR(3 downto 0);
            A, B : in STD_LOGIC_VECTOR(15 downto 0);
            result : out STD_LOGIC_VECTOR(15 downto 0);
            carry, zero, negative, overflow : out STD_LOGIC);
end alu;

architecture alu_one of alu is
    signal value : STD_LOGIC_VECTOR(16 downto 0) := "00000000000000000";
    signal useflag : STD_LOGIC := '0';

begin
    process(A, B, op) begin
        case op is
            when "0001" => value <= '0' & B; --databus
                           useflag <= '1';
            when "0011" => value <= "00000000000000000"; --nollställ
                           useflag <= '1';
            when "0100" => value <= STD_LOGIC_VECTOR('0' & unsigned(A) + unsigned(B)); --add
                           useflag <= '1';
            when "0101" => value <= ('0' & A) - B; --sub
                           useflag <= '1';
            when "0110" => value <= '0' & A and '0' & B; -- and
                           useflag <= '1';
            when "0111" => value <= '0' & A or '0' & B; -- or
                           useflag <= '1';
            when "1000" => value <= STD_LOGIC_VECTOR('0' & unsigned(A) + unsigned(B)); --add noflag
                           useflag <= '0';
            when "1001" => value <= a & '0'; -- ASL/LSL
                           useflag <= '1';
            when "1011" => value <= a(0) & a(15) & a(15 downto 1); -- ASR
                           useflag <= '1';
            when "1101" => value <= a(0) & '0' & a(15 downto 1); -- LSR
                           useflag <= '1';
            when others => value <= '0' & A; -- AR
                           useflag <= '0';
        end case;
    end process;
    
    process(clk) begin
    --process(value, useflag) begin
        if rising_edge(clk) then
            result <= value(15 downto 0);
            if useflag = '1' then
                if value(15 downto 0) = X"0000" then
                    zero <= '1';
                else
                    zero <= '0';
                end if;
                if value(16) = '1' then carry <= '1';
                else carry <= '0'; 
                end if;
                if value(15) = '1' then negative <= '1'; 
                else negative <= '0'; 
                end if;
                if value(16) /= value(15) then overflow <= '1';
                else overflow <= '0';
                end if;
            end if; 
        end if;
    end process;
end alu_one;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity cpu is
    Port (clk,rst : in  STD_LOGIC;
        sw: in STD_LOGIC_VECTOR(7 downto 0);
        seg: out  STD_LOGIC_VECTOR(7 downto 0);
        an : out  STD_LOGIC_VECTOR (3 downto 0);
        led : out STD_LOGIC_VECTOR (7 downto 0);
        vr_we : out STD_LOGIC;
        vr_addr : out STD_LOGIC_VECTOR(4 downto 0);
        vr_i : out STD_LOGIC_VECTOR(15 downto 0);
        vr_o : in STD_LOGIC_VECTOR(15 downto 0);
        fV: in STD_LOGIC;
        up, right, down, left : in STD_LOGIC);
end cpu;

architecture cpu_one of cpu is

    component leddriver
        Port ( clk,rst : in  STD_LOGIC;
           seg : out  STD_LOGIC_VECTOR(7 downto 0);
           an : out  STD_LOGIC_VECTOR (3 downto 0);
           led : out STD_LOGIC_VECTOR (7 downto 0);
           value : in  STD_LOGIC_VECTOR (15 downto 0);
           ledval : in STD_LOGIC_VECTOR (7 downto 0));
    end component;

    component alu
        Port (clk : in STD_LOGIC;
            op : in STD_LOGIC_VECTOR(3 downto 0);
            A, B : in STD_LOGIC_VECTOR(15 downto 0);
            result : out STD_LOGIC_VECTOR(15 downto 0);
            carry, zero, negative, overflow : out STD_LOGIC);
    end component;

    signal databus : STD_LOGIC_VECTOR(15 downto 0) := X"0000";

    -- Registers
    signal rASR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rIR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rPC : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rDR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rAR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rHR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rSP : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal rLC : STD_LOGIC_VECTOR(7 downto 0) := X"00";

    -- Flags
    signal fZ : STD_LOGIC := '1';
    signal fN : STD_LOGIC := '0';
    signal fC : STD_LOGIC := '0';
    signal fO : STD_LOGIC := '0';
    signal fL : STD_LOGIC := '0';

    -- Primary memory
    type PrimMem_type is array (0 to 2047) of STD_LOGIC_VECTOR(15 downto 0);
    signal PrimMem : PrimMem_type := (  0=> X"0100",1=> X"0000",2=> X"0110",3=> X"00d0",4=> X"0120",5=> X"0001",6=> X"0130",7=> X"0002",8=> X"0510",9=> X"0020",10=> X"0510",11=> X"0021",12=> X"0500",13=> X"0022",14=> X"0500",15=> X"0023",16=> X"0500",17=> X"0024",18=> X"0500",19=> X"0025",20=> X"0500",21=> X"0026",22=> X"0500",23=> X"002b",24=> X"0500",25=> X"002c",26=> X"0520",27=> X"002d",28=> X"0530",29=> X"002e",30=> X"0d00",31=> X"0037",32=> X"0000",33=> X"0000",34=> X"0000",35=> X"0000",36=> X"0000",37=> X"0000",38=> X"0000",39=> X"0000",40=> X"0000",41=> X"0000",42=> X"0000",43=> X"0000",44=> X"0000",45=> X"0000",46=> X"0000",47=> X"0000",48=> X"0000",49=> X"0000",50=> X"0000",51=> X"0000",52=> X"0000",53=> X"0000",54=> X"0000",55=> X"3500",56=> X"07ff",57=> X"2500",58=> X"0062",59=> X"2500",60=> X"0073",61=> X"2500",62=> X"00bd",63=> X"2500",64=> X"0106",65=> X"2500",66=> X"014b",67=> X"2500",68=> X"016a",69=> X"2500",70=> X"0189",71=> X"2500",72=> X"01f2",73=> X"2500",74=> X"0267",75=> X"0220",76=> X"002f",77=> X"4120",78=> X"0004",79=> X"0a20",80=> X"0030",81=> X"4120",82=> X"0004",83=> X"0a20",84=> X"0031",85=> X"4120",86=> X"0004",87=> X"0a20",88=> X"0032",89=> X"0230",90=> X"002c",91=> X"0240",92=> X"002b",93=> X"0250",94=> X"0023",95=> X"1c00",96=> X"0d00",97=> X"0039",98=> X"2d00",99=> X"0000",100=> X"0200",101=> X"0035",102=> X"3900",103=> X"0001",104=> X"2100",105=> X"f9c0",106=> X"1900",107=> X"006e",108=> X"0100",109=> X"0280",110=> X"0500",111=> X"0035",112=> X"3100",113=> X"0000",114=> X"2800",115=> X"2d00",116=> X"0000",117=> X"2d10",118=> X"0000",119=> X"0200",120=> X"8000",121=> X"2100",122=> X"0001",123=> X"1900",124=> X"0085",125=> X"0100",126=> X"0020",127=> X"0500",128=> X"0026",129=> X"0100",130=> X"0000",131=> X"0500",132=> X"0025",133=> X"0200",134=> X"8001",135=> X"0210",136=> X"8003",137=> X"2001",138=> X"4d00",139=> X"0098",140=> X"1500",141=> X"00a2",142=> X"0110",143=> X"0002",144=> X"0510",145=> X"002c",146=> X"0110",147=> X"0001",148=> X"0510",149=> X"002b",150=> X"0d00",151=> X"00b8",152=> X"0110",153=> X"0002",154=> X"0510",155=> X"002c",156=> X"0110",157=> X"0000",158=> X"0510",159=> X"002b",160=> X"0d00",161=> X"00b8",162=> X"0210",163=> X"0024",164=> X"2110",165=> X"0000",166=> X"1500",167=> X"00b4",168=> X"5610",169=> X"0023",170=> X"0910",171=> X"0001",172=> X"0510",173=> X"002b",174=> X"0110",175=> X"0001",176=> X"0510",177=> X"002c",178=> X"0d00",179=> X"00b8",180=> X"0110",181=> X"0000",182=> X"0510",183=> X"002c",184=> X"3110",185=> X"0000",186=> X"3100",187=> X"0000",188=> X"2800",189=> X"2d00",190=> X"0000",191=> X"2d10",192=> X"0000",193=> X"0200",194=> X"0023",195=> X"0500",196=> X"0027",197=> X"0200",198=> X"0024",199=> X"0500",200=> X"0028",201=> X"0200",202=> X"0023",203=> X"2200",204=> X"002b",205=> X"1500",206=> X"00d1",207=> X"1900",208=> X"00d9",209=> X"0200",210=> X"0024",211=> X"0a00",212=> X"002c",213=> X"0500",214=> X"0024",215=> X"0d00",216=> X"00ed",217=> X"0200",218=> X"0024",219=> X"3a00",220=> X"002c",221=> X"4d00",222=> X"00e3",223=> X"0500",224=> X"0024",225=> X"0d00",226=> X"00ed",227=> X"5600",228=> X"0024",229=> X"0500",230=> X"0024",231=> X"5600",232=> X"0023",233=> X"0900",234=> X"0001",235=> X"0500",236=> X"0023",237=> X"0200",238=> X"0024",239=> X"2100",240=> X"0018",241=> X"4d00",242=> X"00f7",243=> X"0100",244=> X"0018",245=> X"0500",246=> X"0024",247=> X"0200",248=> X"0024",249=> X"2100",250=> X"000a",251=> X"4d00",252=> X"0101",253=> X"0100",254=> X"0000",255=> X"0500",256=> X"0024",257=> X"3110",258=> X"0000",259=> X"3100",260=> X"0000",261=> X"2800",262=> X"0200",263=> X"0025",264=> X"0500",265=> X"0029",266=> X"0200",267=> X"0026",268=> X"0500",269=> X"002a",270=> X"2d00",271=> X"0000",272=> X"2d10",273=> X"0000",274=> X"0200",275=> X"0025",276=> X"2200",277=> X"002d",278=> X"1500",279=> X"011a",280=> X"1900",281=> X"0122",282=> X"0200",283=> X"0026",284=> X"0a00",285=> X"002e",286=> X"0500",287=> X"0026",288=> X"0d00",289=> X"0136",290=> X"0200",291=> X"0026",292=> X"3a00",293=> X"002e",294=> X"4d00",295=> X"012c",296=> X"0500",297=> X"0026",298=> X"0d00",299=> X"0136",300=> X"5600",301=> X"0026",302=> X"0500",303=> X"0026",304=> X"5600",305=> X"0025",306=> X"0900",307=> X"0001",308=> X"0500",309=> X"0025",310=> X"0200",311=> X"0025",312=> X"2100",313=> X"0001",314=> X"1900",315=> X"0146",316=> X"0200",317=> X"0026",318=> X"2100",319=> X"0008",320=> X"4d00",321=> X"0146",322=> X"0100",323=> X"0008",324=> X"0500",325=> X"0026",326=> X"3110",327=> X"0000",328=> X"3100",329=> X"0000",330=> X"2800",331=> X"2d00",332=> X"0000",333=> X"2d10",334=> X"0000",335=> X"2d80",336=> X"0000",337=> X"0200",338=> X"0024",339=> X"0210",340=> X"0020",341=> X"3d00",342=> X"0003",343=> X"0280",344=> X"0023",345=> X"2180",346=> X"0001",347=> X"1900",348=> X"0160",349=> X"0810",350=> X"0d00",351=> X"0161",352=> X"3810",353=> X"0510",354=> X"0020",355=> X"3180",356=> X"0000",357=> X"3110",358=> X"0000",359=> X"3100",360=> X"0000",361=> X"2800",362=> X"2d00",363=> X"0000",364=> X"2d10",365=> X"0000",366=> X"2d80",367=> X"0000",368=> X"0200",369=> X"0026",370=> X"0210",371=> X"0021",372=> X"3d00",373=> X"0003",374=> X"0280",375=> X"0025",376=> X"2180",377=> X"0001",378=> X"1900",379=> X"017f",380=> X"0810",381=> X"0d00",382=> X"0180",383=> X"3810",384=> X"0510",385=> X"0021",386=> X"3180",387=> X"0000",388=> X"3110",389=> X"0000",390=> X"3100",391=> X"0000",392=> X"2800",393=> X"2d00",394=> X"0000",395=> X"2d10",396=> X"0000",397=> X"2d20",398=> X"0000",399=> X"0200",400=> X"0020",401=> X"0210",402=> X"0021",403=> X"2500",404=> X"01be",405=> X"0500",406=> X"002f",407=> X"0200",408=> X"0020",409=> X"0900",410=> X"000f",411=> X"0210",412=> X"0021",413=> X"2500",414=> X"01be",415=> X"0500",416=> X"0030",417=> X"0200",418=> X"0020",419=> X"0210",420=> X"0021",421=> X"0910",422=> X"000f",423=> X"2500",424=> X"01be",425=> X"0500",426=> X"0031",427=> X"0200",428=> X"0020",429=> X"0900",430=> X"000f",431=> X"0210",432=> X"0021",433=> X"0910",434=> X"000f",435=> X"2500",436=> X"01be",437=> X"0500",438=> X"0032",439=> X"3120",440=> X"0000",441=> X"3110",442=> X"0000",443=> X"3100",444=> X"0000",445=> X"2800",446=> X"2d20",447=> X"0000",448=> X"2d30",449=> X"0000",450=> X"2d40",451=> X"0000",452=> X"2df0",453=> X"0000",454=> X"3d00",455=> X"0004",456=> X"3d10",457=> X"0004",458=> X"0050",459=> X"3d00",460=> X"0004",461=> X"4500",462=> X"0007",463=> X"4110",464=> X"0003",465=> X"0801",466=> X"00f0",467=> X"032f",468=> X"0640",469=> X"0005",470=> X"4500",471=> X"000f",472=> X"0130",473=> X"000f",474=> X"3830",475=> X"0140",476=> X"0001",477=> X"4043",478=> X"4424",479=> X"2120",480=> X"0000",481=> X"1500",482=> X"01e7",483=> X"0100",484=> X"0001",485=> X"0d00",486=> X"01e9",487=> X"0100",488=> X"0000",489=> X"31f0",490=> X"0000",491=> X"3140",492=> X"0000",493=> X"3130",494=> X"0000",495=> X"3120",496=> X"0000",497=> X"2800",498=> X"2d00",499=> X"0000",500=> X"2d10",501=> X"0000",502=> X"2d20",503=> X"0000",504=> X"0200",505=> X"002f",506=> X"2100",507=> X"0001",508=> X"1500",509=> X"0212",510=> X"0200",511=> X"0030",512=> X"2100",513=> X"0001",514=> X"1500",515=> X"0212",516=> X"0200",517=> X"0031",518=> X"2100",519=> X"0001",520=> X"1500",521=> X"0212",522=> X"0200",523=> X"0032",524=> X"2100",525=> X"0001",526=> X"1500",527=> X"0212",528=> X"0d00",529=> X"0260",530=> X"0200",531=> X"002a",532=> X"2200",533=> X"0028",534=> X"4d00",535=> X"021a",536=> X"5100",537=> X"023d",538=> X"0100",539=> X"0000",540=> X"0500",541=> X"0024",542=> X"0210",543=> X"0020",544=> X"4510",545=> X"000f",546=> X"0220",547=> X"0020",548=> X"0200",549=> X"0027",550=> X"2100",551=> X"0001",552=> X"1500",553=> X"0230",554=> X"0130",555=> X"0010",556=> X"3831",557=> X"0823",558=> X"0d00",559=> X"0231",560=> X"3821",561=> X"0520",562=> X"0020",563=> X"0200",564=> X"002a",565=> X"2100",566=> X"0000",567=> X"1500",568=> X"0260",569=> X"0100",570=> X"0000",571=> X"0500",572=> X"0028",573=> X"0100",574=> X"0000",575=> X"0500",576=> X"0026",577=> X"0210",578=> X"0021",579=> X"4510",580=> X"000f",581=> X"0220",582=> X"0021",583=> X"0200",584=> X"0029",585=> X"2100",586=> X"0001",587=> X"1500",588=> X"0253",589=> X"0130",590=> X"0010",591=> X"3831",592=> X"0823",593=> X"0d00",594=> X"0254",595=> X"3821",596=> X"0520",597=> X"0021",598=> X"0100",599=> X"0000",600=> X"0500",601=> X"002a",602=> X"0200",603=> X"0028",604=> X"2100",605=> X"0000",606=> X"1900",607=> X"021a",608=> X"3120",609=> X"0000",610=> X"3110",611=> X"0000",612=> X"3100",613=> X"0000",614=> X"2800",615=> X"2d00",616=> X"0000",617=> X"0200",618=> X"0020",619=> X"0500",620=> X"9000",621=> X"0200",622=> X"0021",623=> X"0500",624=> X"9001",625=> X"0100",626=> X"0002",627=> X"0500",628=> X"9012",629=> X"0100",630=> X"fffd",631=> X"0500",632=> X"9013",633=> X"0200",634=> X"0035",635=> X"0500",636=> X"9014",637=> X"3100",638=> X"0000",639=> X"2800",640=> X"2d00",641=> X"0000",642=> X"0200",643=> X"0021",644=> X"3a00",645=> X"8000",646=> X"0a00",647=> X"8002",648=> X"0500",649=> X"0021",650=> X"0200",651=> X"0020",652=> X"0a00",653=> X"8001",654=> X"3a00",655=> X"8003",656=> X"0500",657=> X"0020",658=> X"3100",659=> X"0000",660=> X"2800",
                                        1600=> X"0006",1601=> X"0000",1602=> X"0020",1603=> X"0000",1604=> X"0000",1605=> X"0000",1606=> X"0000",1607=> X"0000",1608=> X"8006",1609=> X"0000",1610=> X"0020",1611=> X"0000",1612=> X"0000",1613=> X"0000",1614=> X"0000",1615=> X"0000",1616=> X"c03f",1617=> X"f000",1618=> X"0000",1619=> X"0000",1620=> X"0000",1621=> X"0000",1622=> X"0000",1623=> X"0000",1624=> X"c020",1625=> X"0000",1626=> X"0000",1627=> X"0000",1628=> X"0000",1629=> X"0000",1630=> X"0000",1631=> X"0000",1632=> X"fe60",1633=> X"0000",1634=> X"0000",1635=> X"0000",1636=> X"0000",1637=> X"0000",1638=> X"0000",1639=> X"0000",1640=> X"2000",1641=> X"7fdc",1642=> X"03f0",1643=> X"0000",1644=> X"0000",1645=> X"0000",1646=> X"0000",1647=> X"0000",1648=> X"2001",1649=> X"c057",1650=> X"fe18",1651=> X"0000",1652=> X"0000",1653=> X"0000",1654=> X"0000",1655=> X"0000",1656=> X"f9c7",1657=> X"0050",1658=> X"0000",1659=> X"0000",1660=> X"0000",1661=> X"0000",1662=> X"0000",1663=> X"0000",1664=> X"8900",1665=> X"0e50",1666=> X"0000",1667=> X"0000",1668=> X"0000",1669=> X"0000",1670=> X"0000",1671=> X"0000",1672=> X"8900",1673=> X"3a50",1674=> X"0000",1675=> X"0000",1676=> X"0000",1677=> X"0000",1678=> X"0000",1679=> X"0000",1680=> X"89ff",1681=> X"e250",1682=> X"0000",1683=> X"03c0",1684=> X"0000",1685=> X"0000",1686=> X"0000",1687=> X"0000",1688=> X"8000",1689=> X"0250",1690=> X"0000",1691=> X"0f00",1692=> X"0000",1693=> X"0000",1694=> X"0000",1695=> X"0000",1696=> X"8000",1697=> X"0250",1698=> X"0000",1699=> X"3c00",1700=> X"0000",1701=> X"0000",1702=> X"0000",1703=> X"0000",1704=> X"bff8",1705=> X"0250",1706=> X"0318",1707=> X"f000",1708=> X"0000",1709=> X"0000",1710=> X"0000",1711=> X"0000",1712=> X"a008",1713=> X"0240",1714=> X"1fff",1715=> X"c000",1716=> X"0000",1717=> X"0000",1718=> X"0000",1719=> X"0000",1720=> X"afe8",1721=> X"0241",1722=> X"f000",1723=> X"c000",1724=> X"0000",1725=> X"0000",1726=> X"0000",1727=> X"0000",1728=> X"a029",1729=> X"c07f",1730=> X"0000",1731=> X"c000",1732=> X"0000",1733=> X"0000",1734=> X"0000",1735=> X"0000",1736=> X"bff9",1737=> X"7040",1738=> X"0000",1739=> X"c000",1740=> X"0000",1741=> X"0000",1742=> X"0000",1743=> X"0000",1744=> X"8009",1745=> X"1fc0",1746=> X"0000",1747=> X"c000",1748=> X"0000",1749=> X"0000",1750=> X"0000",1751=> X"0000",1752=> X"8009",1753=> X"0040",1754=> X"0000",1755=> X"c000",1756=> X"0000",1757=> X"0000",1758=> X"0000",1759=> X"0000",1760=> X"ff09",1761=> X"0000",1762=> X"0000",1763=> X"c000",1764=> X"0000",1765=> X"0000",1766=> X"0000",1767=> X"0000",1768=> X"0109",1769=> X"0000",1770=> X"0000",1771=> X"c000",1772=> X"0000",1773=> X"0000",1774=> X"0000",1775=> X"0000",1776=> X"0109",1777=> X"0000",1778=> X"0000",1779=> X"c000",1780=> X"0000",1781=> X"0000",1782=> X"0000",1783=> X"0000",1784=> X"0109",1785=> X"000c",1786=> X"0000",1787=> X"0000",1788=> X"0000",1789=> X"0000",1790=> X"0000",1791=> X"0000",1792=> X"0109",1793=> X"0007",1794=> X"0000",1795=> X"0000",1796=> X"0000",1797=> X"0000",1798=> X"0000",1799=> X"0000",1800=> X"0109",1801=> X"0001",1802=> X"ffff",1803=> X"c000",1804=> X"0000",1805=> X"0000",1806=> X"0000",1807=> X"0000",1808=> X"ffc9",1809=> X"3f00",1810=> X"0000",1811=> X"c000",1812=> X"0000",1813=> X"0000",1814=> X"0000",1815=> X"0000",1816=> X"0609",1817=> X"01c0",1818=> X"0000",1819=> X"c000",1820=> X"0000",1821=> X"0000",1822=> X"0000",1823=> X"0000",1824=> X"0609",1825=> X"0070",1826=> X"0000",1827=> X"c000",1828=> X"0000",1829=> X"0000",1830=> X"0000",1831=> X"0000",1832=> X"0609",1833=> X"001f",1834=> X"ff80",1835=> X"c000",1836=> X"0000",1837=> X"0000",1838=> X"0000",1839=> X"0000",1840=> X"0600",1841=> X"0000",1842=> X"00e0",1843=> X"c000",1844=> X"0000",1845=> X"0000",1846=> X"0000",1847=> X"0000",1848=> X"0700",1849=> X"0000",1850=> X"0038",1851=> X"c000",1852=> X"0000",1853=> X"0000",1854=> X"0000",1855=> X"0000",1856=> X"0300",1857=> X"0000",1858=> X"000e",1859=> X"c000",1860=> X"0000",1861=> X"0000",1862=> X"0000",1863=> X"0000",1864=> X"0380",1865=> X"0000",1866=> X"0003",1867=> X"c000",1868=> X"0000",1869=> X"0000",1870=> X"0000",1871=> X"0000",1872=> X"0380",1873=> X"0000",1874=> X"0003",1875=> X"c000",1876=> X"0000",1877=> X"0000",1878=> X"0000",1879=> X"0000",1880=> X"03ff",1881=> X"ff00",1882=> X"0007",1883=> X"c000",1884=> X"0000",1885=> X"0000",1886=> X"0000",1887=> X"0000",1888=> X"0000",1889=> X"01c0",1890=> X"001c",1891=> X"0000",1892=> X"0000",1893=> X"0000",1894=> X"0000",1895=> X"0000",1896=> X"0000",1897=> X"007f",1898=> X"fff0",1899=> X"0000",1900=> X"0000",1901=> X"0000",1902=> X"0000",1903=> X"0000",1904=> X"0000",1905=> X"0000",1906=> X"0000",1907=> X"0000",1908=> X"0000",1909=> X"0000",1910=> X"0000",1911=> X"0000",1912=> X"0000",1913=> X"0000",1914=> X"0000",1915=> X"0000",1916=> X"0000",1917=> X"0000",1918=> X"0000",1919=> X"0000",
                                      others=> X"0000");

    -- Micro memory
    type uMem_type is array (0 to 511) of STD_LOGIC_VECTOR(31 downto 0);
    constant uMem : uMem_type := (  0=>X"04100000",
                                    1=>X"03280000",
                                    2=>X"00000400",
                                    3=>X"0A540200",
                                    4=>X"04180000",
                                    5=>X"03500200",
                                    6=>X"04180000",
                                    7=>X"03100000",
                                    8=>X"03500200",
                                    9=>X"05A00600",
                                    10=>X"05100000",
                                    11=>X"0A300600",
                                    12=>X"15000000",
                                    13=>X"4A000000",
                                    14=>X"07A00600",
                                    15=>X"05400600",
                                    16=>X"00002A0F",
                                    17=>X"00000600",
                                    18=>X"0000220F",
                                    19=>X"00000600",
                                    20=>X"0000240F",
                                    21=>X"00000600",
                                    22=>X"00003816",
                                    23=>X"00000600",
                                    24=>X"1A000000",
                                    25=>X"55000600",
                                    26=>X"09100000",
                                    27=>X"04300000",
                                    28=>X"05420600",
                                    29=>X"00010000",
                                    30=>X"09100000",
                                    31=>X"03400600",
                                    32=>X"09100000",
                                    33=>X"0A320600",
                                    34=>X"00010000",
                                    35=>X"09100000",
                                    36=>X"03A00600",
                                    37=>X"05900600",
                                    38=>X"1A000000",
                                    39=>X"55000000",
                                    40=>X"07A00600",
                                    41=>X"05008000",
                                    42=>X"1A00342D",
                                    43=>X"D0004000",
                                    44=>X"0000322B",
                                    45=>X"07A00600",
                                    46=>X"05008000",
                                    47=>X"1A003432",
                                    48=>X"90004000",
                                    49=>X"00003230",
                                    50=>X"07A00600",
                                    51=>X"15000000",
                                    52=>X"6A000000",
                                    53=>X"07A00600",
                                    54=>X"15000000",
                                    55=>X"7A000000",
                                    56=>X"07A00600",
                                    57=>X"04180000",
                                    58=>X"13000000",
                                    59=>X"4A040000",
                                    60=>X"07100000",
                                    61=>X"03500200",
                                    62=>X"0000260F",
                                    63=>X"00000600",
                                    64=>X"0000280F",
                                    65=>X"00000600",
                                    66=>X"30000000",
                                    67=>X"55000000",
                                    68=>X"07A00600",
                                    69=>X"05008000",
                                    70=>X"00003846",
                                    71=>X"00007246",
                                    72=>X"00000600",
                                    511=>X"00003E00",
                                    others=> X"00000000");

    -- uPC
    signal uPC : STD_LOGIC_VECTOR(8 downto 0) := (others=>'0');
    signal SuPC : STD_LOGIC_VECTOR(8 downto 0) := (others=>'0');

    signal ctrlword : STD_LOGIC_VECTOR(31 downto 0) := X"00000000";
    alias cALU : STD_LOGIC_VECTOR(3 downto 0) is ctrlword(31 downto 28);
    alias cTB : STD_LOGIC_VECTOR(3 downto 0) is ctrlword(27 downto 24);
    alias cFB : STD_LOGIC_VECTOR(3 downto 0) is ctrlword(23 downto 20);
    alias cP : STD_LOGIC is ctrlword(19);
    alias cM : STD_LOGIC is ctrlword(18);
    alias cSP : STD_LOGIC_VECTOR(1 downto 0) is ctrlword(17 downto 16);
    alias cLC : STD_LOGIC_VECTOR(1 downto 0) is ctrlword(15 downto 14);
    alias cSEQ : STD_LOGIC_VECTOR(4 downto 0) is ctrlword(13 downto 9);
    alias cADR : STD_LOGIC_VECTOR(8 downto 0) is ctrlword(8 downto 0);

    type K1_type is array (0 to 63) of STD_LOGIC_VECTOR(8 downto 0);
    signal K1 : K1_type := (0=>"000001001", --MOVE
                            1=>"000001010", --STORE
                            2=>"000001100", --ADD
                            3=>"000001111", --BRA
                            4=>"000010000", --BCS
                            5=>"000010010", --BEQ
                            6=>"000010100", --BNE
                            7=>"000010110", --WVS
                            8=>"000011000", --CMP
                            9=>"000011010", --JSR
                            10=>"000011101", --RTS
                            11=>"000100000", --PUSH
                            12=>"000100010", --POP
                            13=>"000100101", --SSP
                            14=>"000100110", --SUB
                            15=>"000101001", --LSR
                            16=>"000101110", --LSL
                            17=>"000110011", --AND
                            18=>"000110110", --OR
                            19=>"000111110", --BMI
                            20=>"001000000", --BPL
                            21=>"001000010", --INV
                            22=>"001000101", --LWVS  
                            others=>"111111111"); --HULT

    type K2_type is array (0 to 3) of STD_LOGIC_VECTOR(8 downto 0);
    signal K2 : K2_type := (0=>"000000011", --reg-reg
                            1=>"000000100", --imm
                            2=>"000000110", --indir
                            3=>"000111001", --index
                            others=>"000000000");

    type gr_array is array (0 to 15) of STD_LOGIC_VECTOR(15 downto 0);
    signal rGR : gr_array := (others=> X"0000");

    signal tempGR : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal tempPM : STD_LOGIC_VECTOR(15 downto 0) := X"0000";
    signal tempMM : STD_LOGIC_VECTOR(15 downto 0) := X"0000";


    ---------- DEBUG --------
    signal old_step : STD_LOGIC := '0';

begin
    ctrlword <= uMem(conv_integer(uPC));

    led_driver: leddriver port map (clk, rst, seg, an, led, rGR(2), rGR(5)(0) & rGR(4)(0) & "00000" & rGR(3)(0)); --rGR(2) 7-seg, rGR(3) leds
    --led_driver: leddriver port map (clk, rst, seg, an, led, rGR(2), rGR(5)(7 downto 0)); --rGR(2) 7-seg, rGR(3) leds
    alu_instance: alu port map(clk, cALU, rAR, databus, rAR, fC, fZ, fN, fO);
    

    -- *****************************
    -- * CONTROL UNIT              *
    -- *****************************
    process(clk) begin
        if rising_edge(clk) then
            
            -- rst
            if rst = '1' then
                rPC <= X"0000";
                uPC <= "000000000";
            else

                -- LC control
                case cLC is
                    when "01" => rLC <= rLC - 1;
                    when "10" => rLC <= databus(7 downto 0);
                    when "11" => rLC <= cADR(7 downto 0);
                    when others => null;
                end case;

                -- P control
                if cP = '1' then
                    rPC <= rPC + 1; 
                end if;

                -- SP control
                case cSP is
                    when "01" => rSP <= rSP + 1;
                    when "10" => rSP <= rSP - 1;
                    when others => null;
                end case;

                -- SEQ
                case cSEQ is
                    when "00000" => uPC <= uPC + 1;
                    when "00001" => uPC <= K1(conv_integer(rIR(15 downto 10)));
                    when "00010" => uPC <= K2(conv_integer(rIR(9 downto 8)));
                    when "00011" => uPC <= "000000000";
                    when "10000" => uPC <= cADR;
                    when "10001" => if fZ = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10010" => if fZ = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10011" => if fN = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10100" => if fN = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10101" => if fC = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10110" => if fC = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "10111" => if fO = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11000" => if fO = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11001" => if fL = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11010" => if fL = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11011" => if fV = '1' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11100" => if fV = '0' then uPC <= cADR; else uPC <= uPC + 1; end if;
                    when "11101" => 
                        uPC <= cADR; 
                        SuPC <= uPC+1;
                    when "11110" => uPC <= SuPC;
                    when "11111" => null;
                    when others => null;
                end case;
                
                -- FROM BUS
                case cFB is
                    when "0001" => rASR <= databus;
                    when "0010" => rIR <= databus;
                    when "0011" => 
                        if (rASR(15) = '0') then
                            PrimMem(conv_integer(rASR)) <= databus;
                        elsif (rASR(15 downto 12) = X"9") then -- VR
                            vr_i <= databus;
                        end if;
                    when "0100" => rPC <= databus;
                    when "0101" => rDR <= databus;
                    when "0110" => null; -- can't write to uM
                    when "0111" => null; -- can't write to AR
                    when "1000" => rHR <= databus;
                    when "1001" => rSP <= databus;
                    when "1010" => 
                        if cM = '0' then 
                            rGR(conv_integer(rIR(7 downto 4))) <= databus;
                        else
                            rGR(conv_integer(rIR(3 downto 0))) <= databus;
                        end if;
                    when others => null;
                end case;
            end if;
        end if;
    end process;

    with rLC select
    fL <= '0' when X"00",
          '1' when others;

    --process(cFB, rASR, databus) begin
    process(clk) begin
        if rising_edge(clk) then
            if cFB = "0011" and rASR(15 downto 12) = X"9" then -- 9xxx address
                vr_we <= '1';
                --vr_i <= databus;
            else
                vr_we <= '0';
            end if;
        end if;
    end process;

    vr_addr <= rASR(4 downto 0);

    -- TO BUS
    with cTB select
    databus <= rASR when "0001",
                rIR when "0010",
                tempPM when "0011", -- PM/MM
                rPC when "0100",
                rDR when "0101",
                --uMem(conv_integer(uPC)) when "0110",
                rAR when "0111",
                rHR when "1000",
                rSP when "1001",
                tempGR when "1010",
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                --vr_o when "1011",
                X"0000" when others;

    -- PM/MemMap
    with rASR(15) select
    tempPM <= PrimMem(conv_integer(rASR)) when '0',
              tempMM when others;

    -- MemMap
    with rASR select
    tempMM <= "000000000000000" & up when X"8000",
              "000000000000000" & right when X"8001",
              "000000000000000" & down when X"8002",
              "000000000000000" & left when X"8003",
              X"00" & sw when X"8004",
              --X"00" & ledval when X"A000",
              --value when X"A001",
              vr_o when X"9000",vr_o when X"9001",vr_o when X"9002",vr_o when X"9003",
              vr_o when X"9004",vr_o when X"9005",vr_o when X"9006",vr_o when X"9007",
              vr_o when X"9008",vr_o when X"9009",vr_o when X"900A",vr_o when X"900B",
              vr_o when X"900C",vr_o when X"900D",vr_o when X"900E",vr_o when X"900F",
              vr_o when X"9010",vr_o when X"9011",vr_o when X"9012",vr_o when X"9013",
              vr_o when X"9014",vr_o when X"9015",vr_o when X"9016",vr_o when X"9017",
              vr_o when X"9018",vr_o when X"9019",vr_o when X"901A",vr_o when X"901B",
              vr_o when X"901C",vr_o when X"901D",vr_o when X"901E",vr_o when X"901F",
              X"EEEE" when others;

    -- M bit
    with cM select
    tempGR <= rGR(conv_integer(rIR(7 downto 4))) when '0',
              rGR(conv_integer(rIR(3 downto 0))) when others;

end cpu_one;
